    INIT_00 => x"AE544F52030282C7B16E1034E4EDE4AE4B43555404026FC7B16E101FE4EDE4AE",
    INIT_01 => x"4E03020BC8B16EE4AFE4EC62ED62AE544F522D040226C5B16E62AF62ECE4EDE4",
    INIT_02 => x"E4A3104E494D03025FC6B16E84EC3A411F584B43495004021BC8B16E62325049",
    INIT_03 => x"A3104E494D5504061AC6B16E0635D02EE4A31058414D03024DC6B16E0635E02D",
    INIT_04 => x"891F3C3002029DC7B16E0635AE22E4A31058414D5504062CC8B16E0635BF25E4",
    INIT_05 => x"103E300202D6C7B16E5F4FB16E1D530426000083103D3002023EC8B16E891F1D",
    INIT_06 => x"0202E2C7B16E5F4FD927E1A33D0102FBC7B16E891F431D891FB16E0226000083",
    INIT_07 => x"3E55020269C8B16EEE26000083103E3C3003029BC8B16EFFFFCC0327E1A33E3C",
    INIT_08 => x"4FC72DE1A33E010249C8B16E5F4FD422E1A33C5502028AC8B16E5F4FE225E1A3",
    INIT_09 => x"02D2C8B16EE0E4E0A4444E4103020BC9B16E5F4FBA2EE1A33C0102EEC8B16E5F",
    INIT_0a => x"545245564E49060279C8B16EE0E8E0A8524F58030226C9B16EE0EAE0AA524F02",
    INIT_0b => x"A8C8B16EFA261F304958062784300635011F54464948534C060262C5B16E5343",
    INIT_0c => x"45545942080681C9B16EFA261F305644062784300635011F5446494853520602",
    INIT_0d => x"14C7B16E0100832D31020240C9B16E0100C32B310202C4C7B16E891E50415753",
    INIT_0e => x"2D0102B6C9B16EE1E32B010259C9B16E56472F320202BCC8B16E49582A320202",
    INIT_0f => x"19C9B16E4959101F063449580635011F2A3244030267C9B16E0100C35343E1A3",
    INIT_10 => x"B16EE820442F3255440406AFC7B16E101F063456460635011F56472F32440302",
    INIT_11 => x"06D5C9B16EEF2D4D5342410302EDC7B16E0100C3534345544147454E0602ECC9",
    INIT_12 => x"011F1D5F063445544147454E4407029BC9B16EDD2D06354D45544147454E3F07",
    INIT_13 => x"443F080633C9B16EE22D4D53424144040252CAB16EE1A31D00C2101F62ED62A3",
    INIT_14 => x"8900C9101F62ED62E30635011F2B44020216CAB16ECF2D06354D45544147454E",
    INIT_15 => x"C9B16E6632E4A3008200C264EC66ED62A366EC06342D44020201CAB16EE1E300",
    INIT_16 => x"ED3D61E665A616342A4D55030259C8B16E008900C9063562ED62E32B4D0202DE",
    INIT_17 => x"E33D64A6E4A7E4E649008661ED61E33DE4E665A661ED008962EB3D61E664A662",
    INIT_18 => x"626963696469656810008E0634444F4D2F4D5506027DCAB16EE4AF643262AEE4",
    INIT_19 => x"62AE534364ECE2261F306469656962ED0225E4A30620FE1C62EDE4A3082462EC",
    INIT_1a => x"370635FA261F30A0E7062700008C303520364C4C49460402C1C9B16E643264AF",
    INIT_1b => x"C20927A0A080A60F205FE4EDE4AE1062AF1062AE62E33E3C530306C2CAB16E20",
    INIT_1c => x"AF1062AE62E345564F4D430502D4CAB16E30351DED26E4ACB16E303501CA1D00",
    INIT_1d => x"3E45564F4D4306022AC6B16E06353035F826E4ACA0E780E60420E4EDE4AE1062",
    INIT_1e => x"343F31B16E06353035F726E4AC10A2E782E60420AB31E4AE1062AF108B3062AE",
    INIT_1f => x"F8261F30E126A0E1082700008C3035203650494B53040666CBB16E101F203720",
    INIT_20 => x"02FDC8C220F8261F30C627A0E1082700008C303520364E4143530406ABC9DD20",
    INIT_21 => x"4F423E0502DFC8B16E0100C32B52414843050220CCB16E0200C32B4C4C454305",
    INIT_22 => x"00832D5241484305064ACCB16E0200832D4C4C4543050694CBB16E0300C35944",
    INIT_23 => x"74CCB16E4958534C4C454305022ECCB16E0300833E59444F42050690CAB16E01",
    INIT_24 => x"52040266CCB16E0300834B4E494C3E454D414E090423CAB16E53524148430503",
    INIT_25 => x"CBC97EC0DBC7C0CB7ACCAEC9DDC626CCE6C704C64EC80BC7D1C6FFC0BD4C4C4F",
    INIT_26 => x"00DCC2FFC0BD544F4C4C41050258CC7EC0D7C940BCC2A7C4FFC0BD4441500302",
    INIT_27 => x"FFC0BD2C430202EACB7EC04900DCC2B3C52CC6A7C4FFC0BD2C01024CC97EC049",
    INIT_28 => x"CCB16E101F85301FC480E6011F3E454D414E0506A8CA7EC04900F0C21DC6A7C4",
    INIT_29 => x"FFC0BD52454F4421050481CCB16E101FFA2682E460C6011F454D414E3E0506E6",
    INIT_2a => x"040DCDB16E1D5A5801C482E6011F4D4D494004049ECC7EC02CC6AEC913CDD4C3",
    INIT_2b => x"CCB16E1D7EC482E6011F434F5640040460CDB16E891F1D82E6011F3F4D4F4804",
    INIT_2c => x"0405CCB16E1D5A012400C6E1A3E4AFE1A362EC011FE4A34E49485449570602FA",
    INIT_2d => x"BD53433E0304C1CC7EC0E0C937C97CBCC2C4C97ACCFCC397C5FFC0BD50534303",
    INIT_2e => x"00DCC2FFBCC2A1C6A4CDFFC0BD3E5343030482CD7EC03CC6A4CD2F00F0C2FFC0",
    INIT_2f => x"C2DDC6D3CD2F00DCC22ACAD1C6FCC3FFC0BD4B4349502D5343070240CA7EC02F",
    INIT_30 => x"26CE25C300BCC20BC7D1C6FFC0BD4C4C4F522D53430702B9CB7EC0BFCD2F00CB",
    INIT_31 => x"CE7EC0BFCDFBC633CE3DC3BFCD39CE25C300BCC2EAC6D3CDDDC620CE3DC3D3CD",
    INIT_32 => x"38CAF2C738CAF2C7FFC0BD2A4D020237CDB16E891F1D891F0634443E5303020A",
    INIT_33 => x"C775CAD1C6D1C6F2C7FFC0BD4D45522F4D53060252CE7EC086CA50C988C7D8CA",
    INIT_34 => x"4F4D2F4D46060271CD7EC000C848CADDC600C848CA50C90BC7DDC613CB38CA0B",
    INIT_35 => x"9EC850C90BC71FC800C848CA0BC700C813CB38CA0BC775CA10C8D1C6FFC0BD44",
    INIT_36 => x"BD2A01024DCD7EC02BC700C8E0C91FC80BC7B9C9D6CE7BC2F2C72ACAD6CE7BC2",
    INIT_37 => x"020CCB7EC0A1CEDDC646CED1C6FFC0BD444F4D2F040242CE7EC0DBC755CEFFC0",
    INIT_38 => x"2A05029ACE7EC0DBC7F0CEFFC0BD444F4D0302E6CD7EC042C8F0CEFFC0BD2F01",
    INIT_39 => x"7EC042C824CFFFC0BD2F2A02028CCC7EC0A1CEDDC655CED1C6FFC0BD444F4D2F",
    INIT_3a => x"C10DBCC2FFC0BD52430202A0CD7EC03F00F0C2CBC1FFC0BD54494D450402D4CC",
    INIT_3b => x"D6C5FFC0BD4543415053050243CF7EC04100F0C23F00CBC2CCC5CBC10ABCC2CB",
    INIT_3c => x"48CFE6C7A4CF25C300BCC200C8D6C5FFC0BD534543415053060275CF7EC048CF",
    INIT_3d => x"3DC348CFB4C6C2CF25C300BCC2FFC0BD45505954040249CB7EC0DBC79CCF3DC3",
    INIT_3e => x"CBC2CCC53F00CBC2CCC548CF0CBCC2FFC0BD454741500402DDCE7EC0DBC7BACF",
    INIT_3f => x"C1F2C7D6C508BCC2AFC068C4FFC0BD45434150534B434142090634CF7EC04100",
