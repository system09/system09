    INIT_00 => x"0CC2FFC0BD474E49545045434341090434CA7EC03F00DCC2FFBCC2CBC1CBC1CB",
    INIT_01 => x"D4C808BCC27EC0DBC764C73BD07BC2D4C8F2C70DBCC254D07BC228C9D6C5E6C7",
    INIT_02 => x"D07BC2D4C84EC804BCC2F2C7D6C51ED06EC2B9C9F1CF4ED07BC2E6C752D07BC2",
    INIT_03 => x"504543434106026DCE1ED06EC2AEC948CF1DC6D7C975C7E6C71ED06EC2DBC767",
    INIT_04 => x"CB00C8CCC510C8FFC0BD444F4D2F55440606BBCD7EC01BD0CCC500C8FFC0BD54",
    INIT_05 => x"C6D8CAD1C6DBC7D8CA10C8FFC0BD2A55440306E7CF7EC0DDC613CB00C8D1C613",
    INIT_06 => x"0270CA7EC01DC6E0C32B00DCC2FFBCC2FFC0BD444C4F48040222CD7EC0D7C9DD",
    INIT_07 => x"09BCC2E6C7FFC0BD54494749443E0604ABCF7EC02B00CBC2C5CCFFC0BD233C02",
    INIT_08 => x"1FC896D095C6CCC4FFC0BD2301027AD07EC0D7C930BCC2D7C937C907BCC21BC9",
    INIT_09 => x"230202EBCE7EC02FD198C243C954C715D1FFC0BD5323020287CF7EC0CDD0F8D0",
    INIT_0a => x"C2AFC09EC8FFC0BD4E474953040256CF7EC0E0C9F2C7C5CCE0C346C7FFC0BD3E",
    INIT_0b => x"C9CF7EC041D12CD1E3D0FFC0BD474E495254532E55440906F1D07EC0CDD02DBC",
    INIT_0c => x"06AED07EC041D158D11FC82CD1E3D075CA10C8FFC0BD474E495254532E440806",
    INIT_0d => x"D1FFC0BD2E554403068FD07EC0B0CF8ECFE0C95DC854C7FFC0BD455059545205",
    INIT_0e => x"0202CAD17EC0A6D1DDC673D1D1C6FFC0BD522E55440406C8D07EC07BCFB0CF73",
    INIT_0f => x"021ECF7EC0BCD100BCC2FFC0BD2E55020213D17EC07BCFB0CF8AD1FFC0BD2E44",
    INIT_10 => x"D17EC0A6D1DDC68AD1D1C6FFC0BD522E440302A0D17EC0E2D146CEFFC0BD2E01",
    INIT_11 => x"C6FFC0BD522E0202E0D07EC0A6D1DDC673D100BCC2D1C6FFC0BD522E55030229",
    INIT_12 => x"4345440702DFD17EC002D295C6FFC0BD3F010200CF7EC0A6D1DDC68AD146CED1",
    INIT_13 => x"C6CCC410BCC2FFC0BD5845480302B8D17EC02CC6CCC40ABCC2FFC0BD4C414D49",
    INIT_14 => x"554F530602F0D17EC02CC6CCC402BCC2FFC0BD5952414E494206063CCC7EC02C",
    INIT_15 => x"AFE4EC62ED62E3011F474E495254532F070222D27EC043C44EC4FFC0BD454352",
    INIT_16 => x"435441432906049CD2B16E10365E304036284843544143060411D0B16EE1A3E4",
    INIT_17 => x"0469D17EC0E1D270C0CFD2FFC0BD484354414305023ED1B16E5F4F0634443348",
    INIT_18 => x"524F42410502AFD2B16E2037101F4037F926C1A310301F011F574F5248542806",
    INIT_19 => x"6E20C002227AC1062561C1524550505528060473D27EC007D3FFBCC2FFC0BD54",
    INIT_1a => x"AEC91DC6F2C735D389C6E6C764D325C300BCC2FFC0BD524550505505064ED2B1",
    INIT_1b => x"7EC8D1C6E0C954C71FC8FFC0BD455241504D4F43070244D37EC0DBC754D33DC3",
    INIT_1c => x"4F4D0402ECD27EC0AEC9C4C9BFC8AFC0E6C7DDC67EC02BC78CD37BC2C9C76ACB",
    INIT_1d => x"414C50050600D37EC0C0CB7EC09ACBB5D37BC289CD75C7D7C954C7FFC0BD4556",
    INIT_1e => x"A3D2D1C6FFC0BD44524F57040253D17EC0A2D300C834CC1DC654C7FFC0BD4543",
    INIT_1f => x"3CC6B3C454C7E0C9F2C7D1C60ACCDDC600C8F2C7EFCB0BC710C8B7D295C6BFC4",
    INIT_20 => x"BD45535241500502BCD37EC0A7C450C6BFC4E0C9D7C9F2C8E6C7DDC6C2D3A7C4",
    INIT_21 => x"BFC4E0C9D7C9F2C8E6C7DDC6EAC60ACCDDC654C7B7D295C6BFC4A3D2D1C6FFC0",
    INIT_22 => x"C6B16E0635042B5D401F06344B434154533F0606DAD27EC0E0C9F2C7DDC650C6",
    INIT_23 => x"CD49BCC202BCC295C6CCC4FFC0BD455341423F05064DD407D37E1D5C01264DFC",
    INIT_24 => x"D3EABCC292C0D4C8FFC0BD524941503F0506D4D37EC007D3C2BCC264D292C089",
    INIT_25 => x"0802A6D47EC007D3F2BCC292C095C6DAC4FFC0BD504D4F433F0506C8D27EC007",
    INIT_26 => x"4D4F4309046BD37EC04900DCC2B3C52CC6A7C4ACD4FFC0BD2C454C49504D4F43",
    INIT_27 => x"CD7EC02CC6DAC4CCC5FFC0BD5B01030ECF7EC0C8D427C2FFC0BD2928454C4950",
    INIT_28 => x"FFC0BD45524548542D454641530A046CD47EC02CC6DAC4BFC5FFC0BD5D0102CF",
    INIT_29 => x"594C46050400D27EC05CC43D00CBC28BC535D57BC20EC9E0C98BC55CC440BCC2",
    INIT_2a => x"C004D5EAC6DDC64900CBC2E6C73D00CBC2A7C41DD592C095C6DAC4FFC0BD5245",
    INIT_2b => x"FFC0BD2953282204045CD27EC03D00CBC24900CBC25CC4A7C4F4D47EC0E6D4C3",
    INIT_2c => x"C2FFC0BD282E02033CD57EC0B0CF3CC2FFC0BD295328222E050486D27EC03CC2",
    INIT_2d => x"78D57EC0DACCAEC989C6D9D3FFC0BD2C44524F570506BFD47EC0B0CF1FD429BC",
    INIT_2e => x"4F424109049DD37EC0C2D3DACCAEC9F2C7A7C41FD4FFC0BD2C45535241500606",
    INIT_2f => x"06031BD37EC056C207D3FEBCC23100CBC20BC7F8D57BC2FFC0BD295328225452",
    INIT_30 => x"42D5FFC0BD22010739D27EC0C8D522BCC2E6D5E6D442D5FFC0BD2254524F4241",
    INIT_31 => x"42D5FFC0BD222E020319D61ED66EC2FFC0BD225302038FD40FD66EC27DD5E6D4",
    INIT_32 => x"00CBC2E8CCB6C3E8CC00C8A7C4FFC0BD2247534D0406F2D40FD66EC28DD5E6D4",
    INIT_33 => x"0438D67EC0CEC9E0C900C871C504C6FFC0BD48545045440502C1D50FD66EC225",
    INIT_34 => x"45444F4D54494E49080402D57EC089CD8000AFC280BCC2FFC0BD3F5449423805",
    INIT_35 => x"C1BCC2AFC0FFC0BD4C4147454C4C493F0804DCD57EC03300CBC230BCC2FFC0BD",
    INIT_36 => x"BCC2B9C900C83300CBC220BCC2FFC0BD4745525845444E490804AFD67EC007D3",
    INIT_37 => x"BCC2FFC0BD45444F4347455207042ED37EC043C96EC905BCC2B8D60EC9F2C703",
    INIT_38 => x"4040201006040200535559584442412C107DD5D1C6E0C937C9D6C528C9F2C75A",
    INIT_39 => x"45444F4D2B0504DCD407D3C1BCC27EC089C6D7C932D77BC20ACCDDC610C8CEC9",
    INIT_3a => x"040ED27EC037C90FBCC292C0E2C850BCC237C9F000AFC2E6C7D7C918C4FFC0BD",
    INIT_3b => x"AFC200C88AD77BC286D6E6C7E0C9D7C902BCC2A7C400C8FFC0BD4C4552435005",
    INIT_3c => x"C0BD544553464F43060497D67EC0E8CCFDCC00C8B9C97EC0FDCCFDCC37C9FE00",
    INIT_3d => x"10BCC2F0BCC2F2C77EC0DBC7FDCC43C904BCC237C9F000AFC2B8D798C2F2C7FF",
    INIT_3e => x"CC43C937C91FBCC200C837C960BCC2E3D77BC237C9ABC837C910BCC2F2C789CD",
    INIT_3f => x"04FFD57EC0E8CCFDCC7EC0FDCCFDCC37C9FE00AFC2F7D77BC286D6F2C77EC0FD",
