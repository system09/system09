    INIT_00 => x"0816E02F3DC1BD3F3E02087EDF2C3DC1BD3F3C020804DF2A3DC1BD3F3C300308",
    INIT_01 => x"DD013DC1BD58010894DF003DC1BD44010820E07EC050C901BCC2FFC0BD4F4E02",
    INIT_02 => x"43500208B1DD043DC1BD530108E1DF033DC1BD550108ECDF023DC1BD59010827",
    INIT_03 => x"3DC1BD52434303084BE0093DC1BD42010801E0083DC1BD410108D6DF053DC1BD",
    INIT_04 => x"8118DABD2B2B290308AFDE8018DABD2B29020867E00B3DC1BD5044020839E00A",
    INIT_05 => x"30E08418DABD29010842E08318DABD292D2D030898E08218DABD292D02088EE0",
    INIT_06 => x"0C040CE08B18DABD294402085DE08618DABD2941020879E08518DABD29420208",
    INIT_07 => x"023CDF7EC02029028DD5C3C02820028DD5FFC0BD455A49534548544E45524150",
    INIT_08 => x"12E198C2E6C7B9C902D24EC8E6C76ED6AFC06ED67BCFECE054D4FFC0BD532E02",
    INIT_09 => x"F3D14EC8E6C76ED6AFC06ED67BCFECE054D4FFC0BD532E550306B8E07EC0DBC7",
    INIT_0a => x"7BC20EC9F2C7FDBCC2FFC0BD47534D2E040600E17EC0DBC73AE198C2E6C7B9C9",
    INIT_0b => x"7BC295C6E6C795C626CC7AE16EC2B6C37EC0B0CFB4C60BC47BCFAFC0AEC970E1",
    INIT_0c => x"73654D0A8DD5ECE0AFC0C9C7B0CFB4C626CC26CC76E17BC2D4C895C654C78CE1",
    INIT_0d => x"BCC28DC454D472D4FFC0BD4B4F2E0304F6DF7EC03CD200BCC220232065676173",
    INIT_0e => x"CF4B4F20038DD5DFE16EC26B6F20038DD5D9E17BC295C6DAC4DFE17BC237C901",
    INIT_0f => x"C42BE1FFE17BC237C904BCC28DC4FFE16EC203E1F2E17BC237C902BCC28DC459",
    INIT_10 => x"3CD200BCC264D2E6C795C6CCC492C0D4C895C6CCC40ABCC2AFC037C908BCC28D",
    INIT_11 => x"C53B00CBC2E6C766C5FFC0BD59524555510502A3E07EC02029028DD52CC6CCC4",
    INIT_12 => x"C5FFC0BD4C4C49464552060270E07EC07BCF2CC6BFC400BCC23900CBC281D0A7",
    INIT_13 => x"C0BD3E44524F57050627E17EC0CCC57EC0BFC534E2B5E171E27BC2D4C84EC466",
    INIT_14 => x"07D3F0BCC2A0E298C25CE2D1C6DBC77EC042C891E27BC289C6E6C7D9D3E6C7FF",
    INIT_15 => x"CB580FC401E85886E858891F84A6011F4441455248540604B1E181E26EC2DDC6",
    INIT_16 => x"54C75DC820BCC2AEC989C6E6C7FFC0BD454D414E444E4946080484E0B16E1D03",
    INIT_17 => x"42C8EAE298C26ACB75C7E6C7FEE27BC2E6C795C696CCECE26EC2B0E2F2C74AD3",
    INIT_18 => x"C200C8CCC563E37BC2E6C7EAC6FFC0BD44524F57444E49460804D5E07EC042C8",
    INIT_19 => x"E37BC2D1C6E0C9F2C7DDC642C80ACC76CD42C875C718C795C650CC96CC29E36E",
    INIT_1a => x"C813CDE6C742C863E37BC2E6C7DBC723E398C237C90BC765CDE6C7E6C742C845",
    INIT_1b => x"F2C75BC5F0C3AFC0E6C7D0E2E6C7FFC0BD444E4946040207E37EC039C752CD00",
    INIT_1c => x"A7C4D1C6FFC0BD5453494C44524F572D4843524145530F022EE27EC010E3E0C9",
    INIT_1d => x"C0E6C710E301BCC21DC610C813CDA7C4C3E37BC2F2C7DDC6D0E2E6C7A7C4C2D3",
    INIT_1e => x"7EC03500CBC2A7C4FFC0BD4E4F495443455321080465DE7EC042C8DBC7CCC592",
    INIT_1f => x"E8CCAFC2E6D404E47BC289CD80BCC28000AFC2E6C7FFC0BD2C54494C0404A9E2",
    INIT_20 => x"95C6DAC4FFC0BD4C41524554494C0703C1E07EC0D5E3FDCCBCC2E6D47EC0D5E3",
    INIT_21 => x"E3E8E300C8AFC095C6DAC4FFC0BD4C41524554494C320803DFE07EC0E8E3AFC0",
    INIT_22 => x"FFC0BD3E544947494406064FE17EC04500CBC2FFC0BD4B4F3E0306E3E37EC0E8",
    INIT_23 => x"C296E47BC20EC9F2C710BCC284E47BC20EC9F2C709BCC2E0C930BCC20BC7D1C6",
    INIT_24 => x"B5DF7EC0CCC5DDC6DBC77EC02BC7BFC596E47BC20EC995C6CCC4E6C7E0C907BC",
    INIT_25 => x"CCC488C7D1C6D3E47BC25DE489C6F2C7AFC0E6C7FFC0BD5245424D554E3E0702",
    INIT_26 => x"53554E494D0B0478E27EC0DBC7ACE46EC2B7D201BCC288C7C5CADDC6B2D095C6",
    INIT_27 => x"D201BCC205E57BC2D4C82DBCC289C6F2C705E57BC2E6C7FFC0BD3F4E4749532D",
    INIT_28 => x"88C7E6C7CCC5FFC0BD5245424D554E544F443E0A0455E27EC0CCC57EC0BFC5B7",
    INIT_29 => x"00CBC2E6C7A9E4AEC992C046CE43C9D4C82EBCC289C6F2C733E598C2E6C7B9C9",
    INIT_2a => x"E47EC0A9E4B7D201BCC24700CBC2E6C792C0E2C82EBCC289C6F2C7AFC0E6C747",
    INIT_2b => x"7EC02BC7CCC580E57BC242C817E5D1C6E6E4FFC0BD3F5245424D554E44080629",
    INIT_2c => x"C995C6DAC4AFE57BC2C9C76FE3FFC0BD4C4156450404CCE37EC0BFC586CADDC6",
    INIT_2d => x"E57BC29AC4CBE57BC26BE5A1C6B3C4DBC77EC070C07EC0E8CCABE57BC29EC837",
    INIT_2e => x"71C5FFC0BD504F4F4C2D4B4F0704ADE007D3C3BCC27EC019E4DBC77EC032E4C5",
    INIT_2f => x"D4F8C5FFC0BD544955510402A3DEE8E56EC290E57EE2D6C52CC650CC50CC7CC5",
    INIT_30 => x"CF54E17BCFB0CFA1C6B3C41DE698C260C9E6C7A0D659CFF2D2DBE5AFC234E2F4",
    INIT_31 => x"0526C8FF8310B16E0635042600008310574F52485405026AE3FFE56EC2E5C57B",
    INIT_32 => x"3B00CBC23900CBC2FFC0BD544552505245544E49090496DE07D37EFAE57E0635",
    INIT_33 => x"02DAE47EC0DBC76BE698C289C6E6C7D9D3D6C590E56DE66EC22CC6BFC400BCC2",
    INIT_34 => x"BFC4DDC6F2D255E6AFC2D1C695C6BFC4EAC6A3D2FFC0BD455441554C41564508",
    INIT_35 => x"C292C0FFC0BD444E554F463F060480E67EC030E63B00CBC23900CBC2FBC62CC6",
    INIT_36 => x"C0BD52414843040289E37EC0BAE66FE37EE2D6C5FFC0BD2701028BE507D3F3BC",
    INIT_37 => x"CBE07EC019E4DEE6FFC0BD5D524148435B0603F5E57EC089C6AEC97EE2D6C5FF",
    INIT_38 => x"D429BCC2FFC0BD280103C7E27EC019E437C91FBCC2DEE6FFC0BD4C5254430407",
    INIT_39 => x"29BCC289C6B9C9D7C9A3D244E77BC295C6BFC492C00EC943C495C6BFC446C71F",
    INIT_3a => x"060254E07EC02CC6BFC443C4FFC0BD5C010356E47EC01CE798C25CE292C0D4C8",
    INIT_3b => x"26CC80E77BC20BC703BCC2A7C4D1C6E6C7D0E27EE2D6C5FFC0BD455441455243",
    INIT_3c => x"65520B8DD559CFB7E77BC2DDC600BCC22CC6C0CBAEC989C6F2C7A7C4E6C7DACC",
    INIT_3d => x"C7A7C41DC6B9C9A7C443C98000AFC27BCFB0CFB4C6A7C420676E696E69666564",
    INIT_3e => x"C989C6F2C789C65BC5B9C9A7C42CC600C8A7C42CC696CCA7C495C6E6C7B0E2E6",
    INIT_3f => x"4304045FE77EC0D5E311C16ADBCCC5DACCAEC989C62900CBC2A7C41DC600C843",
