--*******************************************************
--
-- NOICE09 Monitor ROM for the 6809
-- noice09_rom2k_b4.vhd
-- John Kent
-- 4th July 2006
--
--*******************************************************
--
-- Using 4 x RAMB4_S8 found in the XC2S300e
-- NOICE09 assumes an ACIA at $E000
-- and Monitor RAM from $F000 to $F7FF
-- The monitor starts at $FC00
-- The first 1K of ROM is empty and may
-- be used for other purposes
--
-- The Noice monitor has the same entity name
-- as SBUG and KBUG9S so it can be easily exchanged.
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
library unisim;
	use unisim.all;

entity mon_rom is
    Port (
       clk   : in  std_logic;
       rst   : in  std_logic;
       cs    : in  std_logic;
       rw    : in  std_logic;
       addr  : in  std_logic_vector (10 downto 0);
       wdata : in  std_logic_vector (7 downto 0);
       rdata : out std_logic_vector (7 downto 0)
    );
end mon_rom;

architecture rtl of mon_rom is

   signal rdata0 : std_logic_vector (7 downto 0);
   signal rdata1 : std_logic_vector (7 downto 0);
   signal rdata2 : std_logic_vector (7 downto 0);
   signal rdata3 : std_logic_vector (7 downto 0);

   signal ena0 : std_logic;
   signal ena1 : std_logic;
   signal ena2 : std_logic;
   signal ena3 : std_logic;

   signal we : std_logic;

   component RAMB4_S8
    generic (
      INIT_00, INIT_01, INIT_02, INIT_03,
	   INIT_04, INIT_05, INIT_06, INIT_07,
	   INIT_08, INIT_09, INIT_0A, INIT_0B,
      INIT_0C, INIT_0D, INIT_0E, INIT_0F : bit_vector (255 downto 0)
    );

    port (
      clk, we, en, rst : in std_logic;
      addr : in std_logic_vector(8 downto 0);
      di : in std_logic_vector(7 downto 0);
      do : out std_logic_vector(7 downto 0)
    );
  end component RAMB4_S8;

begin

  ROM0 : RAMB4_S8
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0f => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map ( clk => clk,
	            en => ena0,
				   we => we,
				   rst => rst,
				   addr(8 downto 0) => addr(8 downto 0),
               di(7 downto 0)   => wdata,
				   do(7 downto 0)   => rdata0(7 downto 0)
	);

  ROM1 : RAMB4_S8
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0f => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map ( clk => clk,
	            en => ena1,
				   we => we,
				   rst => rst,
				   addr(8 downto 0) => addr(8 downto 0),
               di(7 downto 0)   => wdata,
				   do(7 downto 0)   => rdata1(7 downto 0)
	);

  ROM2 : RAMB4_S8
    generic map ( 
    INIT_00 => x"ACFC8E1001E07D00E0B7118600E0B70386FA2612121F3000008E20F6CE10321A",
    INIT_01 => x"2AF6B72BF6B72EF6FD0000CC22F6F723F6B710F6CCFA265A81AF1008C600F08E",
    INIT_02 => x"34D1FD7E30F6B7FA862DF6B7828621F6B720F6B724F6FD26F6FD28F6FD2CF6B7",
    INIT_03 => x"FCBD02349035011A903501E0B64FF227018400E0B60D271F308EFCBD00008E10",
    INIT_04 => x"6D20393038363F0100000000008005394C4F3901E0B70235F627028400E0B68E",
    INIT_05 => x"02352AF6B702352BF6B702352DF6B7023520F6B700302E315620726F74696E6F",
    INIT_06 => x"20F6B6103524F6F725F6B7063526F6F727F6B7063528F6F729F6B706352CF6B7",
    INIT_07 => x"25F781F4255FFCBD30F68E20F6CE1037FE7E2EF6F72FF6B7101F1F3002260181",
    INIT_08 => x"FCBDF6265A80A7D8255FFCBD891F0C27008180A7E5228081E9255FFCBD80A7F0",
    INIT_09 => x"812527FD812627FE814227FF8180E680A630F68EC526E0ABB4FEBD0234CE255F",
    INIT_0a => x"FE7E018630F6B7F0861F27F7812027F8812127F9812227FA812327FB812427FC",
    INIT_0b => x"31F68E1091FC8E84FE7E79FE7E4BFE7EF8FD7EE6FD7ED1FD7EA5FD7E8EFD7E92",
    INIT_0c => x"5A80A7A0A6072731F6F703E6021F01E602A69CFE7EF9265AA0A780A6A0E71BC6",
    INIT_0d => x"A63435F9265AA0A780A63434142703C031F6F6021F80A680E680A69CFE7EF926",
    INIT_0e => x"80A7A0A680E731F68E10C620F68E1092FE7E018602200086F7265A0726A0A180",
    INIT_0f => x"041F22F6F623F6B692FE7E4FF9265AA0A780A620F68E100B275D9CFE7EF9265A"
    )
    port map ( clk => clk,
	            en => ena2,
				   we => we,
				   rst => rst,
				   addr(8 downto 0) => addr(8 downto 0),
               di(7 downto 0)   => wdata,
				   do(7 downto 0)   => rdata2(7 downto 0)
	);

  ROM3 : RAMB4_S8
    generic map ( 
    INIT_00 => x"063428F6F629F6B6063426F6F627F6B6063424F6F625F6B606342EF6F62FF6B6",
    INIT_01 => x"1022F6F723F6B7401F3B0234508A2DF6B602342BF6B602342AF6B602342CF6B6",
    INIT_02 => x"A4A6021F01E602A6043420275454C0A7008631F6CED1FD7E21F6B7008620F6CE",
    INIT_03 => x"A6021F84E601A69CFE7EE02631F6F1043031F67CC0A70C260435A4E1A4E703E6",
    INIT_04 => x"40B4FEBD002031F6B7018632F6B792FE7E4FA4A702A6021F84E601A692FE7EA4",
    INIT_05 => x"5A80AB008602CB01E630F68EF1FC7EF8265A7CFCBD80A603CB01E630F68E84A7",
    INIT_06 => x"26508502352BF6B7846E04F0BE0586846E02F0BE0686846E00F0BE078639FB26",
    INIT_07 => x"6E0CF0BE0286846E08F0BE0386846E06F0BE04860234508A04342BF6F67C3409",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000ACFC7E018684",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0f => x"00FCFAFE01FFF3FED8FED1FECAFEC3FE00000000000000000000000000000000"
    )
    port map ( clk => clk,
	            en => ena3,
				   we => we,
				   rst => rst,
				   addr(8 downto 0) => addr(8 downto 0),
               di(7 downto 0)   => wdata,
				   do(7 downto 0)   => rdata3(7 downto 0)
	);

my_noice09_b4 : process ( cs, rw, addr, rdata0, rdata1, rdata2, rdata3 )
begin
		   case addr(10 downto 9) is
			when "00" =>
			   ena0  <= cs;
				ena1  <= '0';
				ena2  <= '0';
				ena3  <= '0';
            rdata <= rdata0;
			when "01" =>
			   ena0  <= '0';
				ena1  <= cs;
				ena2  <= '0';
				ena3  <= '0';
            rdata <= rdata1;
			when "10" =>
			   ena0  <= '0';
				ena1  <= '0';
				ena2  <= cs;
				ena3  <= '0';
            rdata <= rdata2;
			when "11" =>
			   ena0  <= '0';
				ena1  <= '0';
				ena2  <= '0';
				ena3  <= cs;
            rdata <= rdata3;
			when others =>
			   null;
			end case;

	 we <= not rw;

end process;

end architecture rtl;

