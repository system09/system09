library IEEE;
   use IEEE.std_logic_1164.all;
   use IEEE.std_logic_arith.all;
library unisim;
   use unisim.vcomponents.all;

entity my_rom is
   port(
      clk      : in  std_logic;
      rst      : in  std_logic;
      cs       : in  std_logic;
      rw       : in  std_logic;
      addr     : in  std_logic_vector(11 downto 0);
      data_in  : in  std_logic_vector(7 downto 0);
      data_out : out std_logic_vector(7 downto 0)
   );
end my_rom;

architecture rtl of my_rom is
   type d_type is array( 0 to 1 ) of std_logic_vector(7 downto 0);
   type p_type is array( 0 to 1 ) of std_logic_vector(0 downto 0);
   signal do : d_type;
   signal dp : p_type;
   signal en : std_logic_vector(1 downto 0);
   signal we : std_logic;
begin
   ROM0: RAMB16_S9
      generic map (
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0f => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1f => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2f => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3f => x"0000000000000000000000000000000000000000000000000000000000000000",
      )
      port map (
         do      => do(0),
         dop     => dp(0),
         addr    => addr(10 downto 0),
         clk     => clk,
         di      => data_in,
         dip     => dp(0),
         en      => en(0),
         ssr     => rst,
         we      => we
      );
   ROM1: RAMB16_S9
      generic map (
    INIT_00 => x"A780A610C6C0DF8E105FFE8E2EFA17FB1BFB8CFBCBFCB6FC98FC9EFC61F814F8",
    INIT_01 => x"17431FE4A7D0866AAFDD8C30FB265AE26F0CC65B0117E0DFBF00E08EF9265AA0",
    INIT_02 => x"031792FE8E090417F62A5A19048B0327856D0DC64FD0DF8E4403176FFE8EA004",
    INIT_03 => x"17408B981F5004175E86092C2081891FF1270D817F84340417B0021799FE8E2B",
    INIT_04 => x"20ED02179BFE8EF5265FFE8C02300F2780E126FE8E20C0022F60C14404174904",
    INIT_05 => x"17A4A60C0417A20317211F620217A1FE8E121F2D296803173B341FBC2094ADC0",
    INIT_06 => x"27A4A1A4A7390F260D8117275E81DD271881E127088111285B0317040417A203",
    INIT_07 => x"08031705201F30C0DF8E321F9F0217BE203F31C2202131E203173F86E5031708",
    INIT_08 => x"279703170527E4AC011FF0C4201F0634F0C41000C3101F390124E1AC20340629",
    INIT_09 => x"265A8B031729031780A610C69303172B0317E4AEEB0117A1FE8E103439623203",
    INIT_0a => x"29B40217BC20EE265A7403172E8602237E810425208180A610C6E1AE830317F5",
    INIT_0b => x"3984A73F86A4AFA0A709273F8184A60F271035558DFFFF8E10341A24C0DF8C1E",
    INIT_0c => x"4AAF0427268D1F304AAE431F39FB265A188D08C6E3DF8E104303163F86460317",
    INIT_0d => x"A7A0A7A0A7FF8684A7A4A604263F8184A60A24C0DF8C21AEB9FE16450217068D",
    INIT_0e => x"0186398D46E0B7E086408D393D3139F7265A0427A1ACA0A608C6E3DF8E1039A0",
    INIT_0f => x"178D47E0B7208645E0B744E0B743E0B74F42E0B701862D8D47E0B7EF8641E0B7",
    INIT_10 => x"E0B6F926808547E0B63B341F4AAF00C08EF42600C28C80A740E0B6218D00C08E",
    INIT_11 => x"54545454A6E6D0DF8E104444444462A6363439F927088547E0B639F227408547",
    INIT_12 => x"11868435FD265A20C60434B63562E762EA62A70F8462A65858585853A6E6E4E7",
    INIT_13 => x"1726290234A80117F12631813D273981230217F92653812A0217E2DF7F680217",
    INIT_14 => x"27E46AE0EB02340C2904358E01170434E46AE46AE4EBE0EBE0E6103421299101",
    INIT_15 => x"30344A0117E26F1202161386E2DF731A02173F86BA27FFC102355FEB2080A705",
    INIT_16 => x"20C6022320008310062762A3E4ECF901171286E4FCBDE4AF0130492562AC4D29",
    INIT_17 => x"6A65011780A684EB63EB62EB68011762AE750117981F03CB2F0017E2FE8E64E7",
    INIT_18 => x"93FE8E10347120028D396532B701171486C326E4AC62AF5B0117981F53F52664",
    INIT_19 => x"EB8DE78D618D394AAF0229F68DF28D910017E50016F80016A101169035690017",
    INIT_1a => x"8DC68D498D3944AF0229D58DD18D5E8D3946AF0229E08DDC8D728D3948AF0229",
    INIT_1b => x"A58D5F8D3941A70229B18DB08D588D3942A70229BC8DBB8D6C8D3943A70229C7",
    INIT_1c => x"B1FE8EBF0016311FF48DA5FE8E39F726048180A63F011739C4A7808A0429A68D",
    INIT_1d => x"46AECE8DB7FE8EE12044AED78DBDFE8EB4001643A6E18DC3FE8EF42048AEEA8D",
    INIT_1e => x"D3FE8ED02042A6B38DCEFE8ED92041A6BC8DC9FE8ECF204AAEC58DABFE8ED820",
    INIT_1f => x"17FF17A1FE8EBF8DB88DB08DA98DA18D27FF17A1FE8E900016DAFE8EC4A6AA8D",
    INIT_20 => x"A710343C29088D011F42290E8DB800172D86121F4D29098DD520CE8DC78DC08D",
    INIT_21 => x"032239811D2530815B8D39E0AB04342829078D891F484848483229118D903561",
    INIT_22 => x"0235103439021A39578003226681072561813937800322468112254181393080",
    INIT_23 => x"80A608C602345120078B022F3981308B0F840235048D4444444402340235028D",
    INIT_24 => x"10342D207F84048D0627E2DF7D00F09F6E8235F1265A3F8D438D2D860225E468",
    INIT_25 => x"05260185E0DF9FA60234903501A6EE27018584A620E08E0926018584A6E0DFBE",
    INIT_26 => x"01A70235F6260885FA27028584A6E0DFBE1234498D2086008D8235018520E0B6",
    INIT_27 => x"FBDFFD0000CC30E08E39E2DFB7FF86016D84A7118684A70386E0DFBE138D9035",
    INIT_28 => x"0427FEDF7D30E08E16345986028D1B86FEDF7F01E702C6FDDFFD04E703E702A7",
    INIT_29 => x"0027101A815A271B81342708819635AF001784A70520098D042420810D20608D",
    INIT_2a => x"16792619C15CFBDFFC45260A810F270B8124270C81890027100D81382716817C",
    INIT_2b => x"0000CC5820212750814CFBDFB662204A2C27FBDFB66D205A34275DFBDFFC8F00",
    INIT_2c => x"FDDF7D39FEDF7F39FEDFB704263D81312754816E27598114273DC1FEDFF65620",
    INIT_2d => x"0000CC1B20E12218C120C0FDDF7FFDDFF6ED224F812080FEDF7F39FDDFB70426",
    INIT_2e => x"3903E702A7FBDFFDFCDFF64F39FEDF7FF726508102A74C84E720C6FBDFB6168D",
    INIT_2f => x"2086FBDFF604E75F012519C15C04E6E78D5AEA2619C15C4FF02650814CFBDFFC",
    INIT_30 => x"FBDFF75FE4205F03E7FCDFF7082719C15CFCDFF6F42650C15C84A702E7FBDFF7",
    INIT_31 => x"F94245FB1950FB183AFB152EFB105BFB047CFB0366FB0271FB0139FEDFF702E7",
    INIT_32 => x"F98FFC55D5F94488F958F1F853EAFB52A8F84DB9FA505EFA4CA5F847FDF8455C",
    INIT_33 => x"382E312047554239305359530000000A0DFFFFFFFF94F9A7F8A7F8A7F8A7F894",
    INIT_34 => x"3F54414857043E040000000A0D4B04202D2052455452415453335320524F4620",
    INIT_35 => x"492020043D59492020043D53552020043D43502020043D5053202004202D2004",
    INIT_36 => x"5A4E4948464504203A43432020043D422020043D412020043D50442020043D58",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000431534356",
    INIT_38 => x"300B2784AC1084AF1084EEAA558E10A0D08E84A7F086FB264A80A70F86F0FF8E",
    INIT_39 => x"2DA7D0DF8E10C0DFCE10FDFFB74444444443101F84EFD620ED26A0F08C00F089",
    INIT_3a => x"1084AF10AA558E1084EE2227A0F08C00F08930FB2A4AA66F0C862FA7F0862E6F",
    INIT_3b => x"2EA7D0DF8E10F186D520A5A70F88891F44444444101FD0DF8E1084EFE92684AC",
    INIT_3c => x"8EF32D0C814C80E7A66F0427A6E6211F4F2CE7A66F1420F92A4A0526A6E60C86",
    INIT_3d => x"9F6EC6DF9F6EC4DF9F6EC0DF9F6E62F816E2DFF753F9265A80A7A0A610C6F0FF",
    INIT_3e => x"0822CEDFBC8B300F27FFFF8CCCDFBE49584F4AAF80E64AAE431FCADF9F6EC8DF",
    INIT_3f => x"00FFB2FFC2FFBEFFBAFFB6FFC6FFB2FFC2DF9F6E42EE1F37F16E44AEC4EC1034"
      )
      port map (
         do      => do(1),
         dop     => dp(1),
         addr    => addr(10 downto 0),
         clk     => clk,
         di      => data_in,
         dip     => dp(1),
         en      => en(1),
         ssr     => rst,
         we      => we
      );
   rom_decode: process(rw, addr, do)
   begin
      we <= not rw;
      en <= (others => '0');
      case( addr(11 downto 11)) is
      when "0" =>
          en(0)   <= cs;
          data_out <= do(0);
      when "1" =>
          en(1)   <= cs;
          data_out <= do(1);
      when others =>
          data_out <= (others=>'0');
      end case;
   end process;
end architecture rtl;

