library IEEE;
   use IEEE.std_logic_1164.all;
   use IEEE.std_logic_arith.all;
library unisim;
   use unisim.vcomponents.all;

entity SYS09BUG_F000 is
   port(
      clk    : in  std_logic;
      rst    : in  std_logic;
      cs     : in  std_logic;
      rw     : in  std_logic;
      addr   : in  std_logic_vector(10 downto 0);
      rdata  : out std_logic_vector(7 downto 0);
      wdata  : in  std_logic_vector(7 downto 0)
   );
end SYS09BUG_F000;

architecture rtl of SYS09BUG_F000 is

   type data_array is array(0 to 3) of std_logic_vector(7 downto 0);
   signal xdata : data_array;
   signal en : std_logic_vector(3 downto 0);
   signal we : std_logic;

component RAMB4_S8
generic (
   INIT_00, INIT_01, INIT_02, INIT_03,
   INIT_04, INIT_05, INIT_06, INIT_07,
   INIT_08, INIT_09, INIT_0A, INIT_0B,
   INIT_0C, INIT_0D, INIT_0E, INIT_0F : bit_vector (255 downto 0)
    );
   port (
      clk, we, en, rst : in std_logic;
      addr : in std_logic_vector(8 downto 0);
      di   : in std_logic_vector(7 downto 0);
      do   : out std_logic_vector(7 downto 0)
      );
     end component RAMB4_S8;

   begin

   ROM00: RAMB4_S8
      generic map (
         INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0a => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0b => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0c => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0d => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0e => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0f => x"0000000000000000000000000000000000000000000000000000000000000000"
      )
      port map (
         clk     => clk,
         en      => en(0),
         we      => we,
         rst     => rst,
         addr    => addr(8 downto 0),
         di      => wdata,
         do      => xdata(0)
      );

   ROM01: RAMB4_S8
      generic map (
         INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0a => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0b => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0c => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0d => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0e => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0f => x"0000000000000000000000000000000000000000000000000000000000000000"
      )
      port map (
         clk     => clk,
         en      => en(1),
         we      => we,
         rst     => rst,
         addr    => addr(8 downto 0),
         di      => wdata,
         do      => xdata(1)
      );

   ROM02: RAMB4_S8
      generic map (
         INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0a => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0b => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0c => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0d => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0e => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0f => x"0000000000000000000000000000000000000000000000000000000000000000"
      )
      port map (
         clk     => clk,
         en      => en(2),
         we      => we,
         rst     => rst,
         addr    => addr(8 downto 0),
         di      => wdata,
         do      => xdata(2)
      );

   ROM03: RAMB4_S8
      generic map (
         INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0a => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0b => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0c => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0d => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0e => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0f => x"0000000000000000000000000000000000000000000000000000000000000000"
      )
      port map (
         clk     => clk,
         en      => en(3),
         we      => we,
         rst     => rst,
         addr    => addr(8 downto 0),
         di      => wdata,
         do      => xdata(3)
      );

   rom_glue: process (cs, rw, addr, xdata)
   begin
      en <= (others=>'0');
      case addr(10 downto 9) is
      when "00" =>
         en(0)  <= cs;
         rdata  <= xdata(0);
      when "01" =>
         en(1)  <= cs;
         rdata  <= xdata(1);
      when "10" =>
         en(2)  <= cs;
         rdata  <= xdata(2);
      when "11" =>
         en(3)  <= cs;
         rdata  <= xdata(3);
      when others =>
         null;
      end case;
      we <= not rw;
   end process;
end architecture rtl;

library IEEE;
   use IEEE.std_logic_1164.all;
   use IEEE.std_logic_arith.all;
library unisim;
   use unisim.vcomponents.all;

entity SYS09BUG_F800 is
   port(
      clk    : in  std_logic;
      rst    : in  std_logic;
      cs     : in  std_logic;
      rw     : in  std_logic;
      addr   : in  std_logic_vector(10 downto 0);
      rdata  : out std_logic_vector(7 downto 0);
      wdata  : in  std_logic_vector(7 downto 0)
   );
end SYS09BUG_F800;

architecture rtl of SYS09BUG_F800 is

   type data_array is array(0 to 3) of std_logic_vector(7 downto 0);
   signal xdata : data_array;
   signal en : std_logic_vector(3 downto 0);
   signal we : std_logic;

component RAMB4_S8
generic (
   INIT_00, INIT_01, INIT_02, INIT_03,
   INIT_04, INIT_05, INIT_06, INIT_07,
   INIT_08, INIT_09, INIT_0A, INIT_0B,
   INIT_0C, INIT_0D, INIT_0E, INIT_0F : bit_vector (255 downto 0)
    );
   port (
      clk, we, en, rst : in std_logic;
      addr : in std_logic_vector(8 downto 0);
      di   : in std_logic_vector(7 downto 0);
      do   : out std_logic_vector(7 downto 0)
      );
     end component RAMB4_S8;

   begin

   ROM00: RAMB4_S8
      generic map (
         INIT_00 => x"A780A610C6C07F8E104EFE8ECFFE0DFB11FB82FBBDFCA8FC8AFC90FC4BF814F8",
         INIT_01 => x"17431FE4A7D0866AAFDD8C30FB265AE26F0CC6450117D07FBF00E08EF9265AA0",
         INIT_02 => x"092C2081891FF1270D817F843C0417BC021783FE8EDE01173A03175EFE8E9204",
         INIT_03 => x"FE8C02300F2780E118FE8E20C0022F60C14C0417510417408B981F5804175E86",
         INIT_04 => x"1F6E02178BFE8E121F2D297403173B341FBC2094ADC020F9021785FE8EF5264E",
         INIT_05 => x"17275E81DD271881E127088111286703170C0417AE0317A4A6140417AE031721",
         INIT_06 => x"321FAB0217BE203F31C2202131EA03173F86ED03170827A4A1A4A7390F260D81",
         INIT_07 => x"F0C4201F0634F0C41000C3101F390124E1AC2034062914031705201F30C07F8E",
         INIT_08 => x"10C69B0317370317E4AEF701178BFE8E103439623203279F03170527E4AC011F",
         INIT_09 => x"03172E8602237E810425208180A610C6E1AE8B0317F5265A93031735031780A6",
         INIT_0a => x"273F8184A60F2710355B8DFFFF8E10341A24C07F8C1E29C00217BC20EE265A7C",
         INIT_0b => x"431F39FB265A1E8D08C6D37F8E104B03163F864E03173984A73F86A4AFA0A709",
         INIT_0c => x"A60A24C07F8C21AEB3FE16ED7FBF00008E5102170C8D4AAF04272C8D1F304AAE",
         INIT_0d => x"265A0427A1ACA0A608C6D37F8E1039A0A7A0A7A0A7FF8684A7A4A604263F8184",
         INIT_0e => x"7FBFE7F98EEB7FBFC07FBEED7FBF1429390217EE02171C295F0117393D3139F7",
         INIT_0f => x"27ED7FBE24273F8184A64AAEEC011770E0B671E0B73686431F392020450017C0"
      )
      port map (
         clk     => clk,
         en      => en(0),
         we      => we,
         rst     => rst,
         addr    => addr(8 downto 0),
         di      => wdata,
         do      => xdata(0)
      );

   ROM01: RAMB4_S8
      generic map (
         INIT_00 => x"3B71E0B73F8673E0B7368670E0B671E0B7368670E0B70D86341FED7FBF1F301F",
         INIT_01 => x"B7368672E0B7008670E0B7FF8673E0B73A8671E0B7328622FE16C07FBFEB7FBE",
         INIT_02 => x"81260217D27F7F6402171186D6FCBD8435FD265A20C604343973E0B73E8671E0",
         INIT_03 => x"E0EBE0E61034212991011726290234A80117F12631813D2739811F0217F92653",
         INIT_04 => x"FFC102355FEB2080A70527E46AE0EB02340C2904358E01170434E46AE46AE4EB",
         INIT_05 => x"E4AF0130492562AC4D2930344A0117E26F0E02161386D27F731602173F86BA27",
         INIT_06 => x"03CB2F0017CCFE8E64E720C6022320008310062762A3E4ECF501171286D6FCBD",
         INIT_07 => x"AF5B0117981F53F526646A65011780A684EB63EB62EB68011762AE750117981F",
         INIT_08 => x"00169D011690356900177DFE8E10347120028D396532B301171486C326E4AC62",
         INIT_09 => x"8DDC8D728D3948AF0229EB8DE78D618D394AAF0229F68DF28D910017E50016F8",
         INIT_0a => x"BB8D6C8D3943A70229C78DC68D498D3944AF0229D58DD18D5E8D3946AF0229E0",
         INIT_0b => x"1739C4A7808A0429A68DA58D5F8D3941A70229B18DB08D588D3942A70229BC8D",
         INIT_0c => x"8DADFE8EF42048AEEA8D9BFE8EBF0016311FF48D8FFE8E39F726048180A63B01",
         INIT_0d => x"204AAEC58D95FE8ED82046AECE8DA1FE8EE12044AED78DA7FE8EB4001643A6E1",
         INIT_0e => x"900016C4FE8EC4A6AA8DBDFE8ED02042A6B38DB8FE8ED92041A6BC8DB3FE8ECF",
         INIT_0f => x"098DD520CE8DC78DC08D17FF178BFE8EBF8DB88DB08DA98DA18D27FF178BFE8E"
      )
      port map (
         clk     => clk,
         en      => en(1),
         we      => we,
         rst     => rst,
         addr    => addr(8 downto 0),
         di      => wdata,
         do      => xdata(1)
      );

   ROM02: RAMB4_S8
      generic map (
         INIT_00 => x"4848483229118D903561A710343C29088D011F42290E8DB400172D86121F4D29",
         INIT_01 => x"22468112254181393080032239811D253081578D39E0AB04342829078D891F48",
         INIT_02 => x"4444444402340235028D0235103439021A395780032266810725618139378003",
         INIT_03 => x"3B8D3F8D2D860225E46880A608C602344D20078B022F3981308B0F840235048D",
         INIT_04 => x"84A620E08E0926018584A6D07FBE10342D207F84048D0627D27F7D8235F1265A",
         INIT_05 => x"34498D2086008D8235018520E0B605260185D07F9FA60234903501A6EE270185",
         INIT_06 => x"A7518684A70386D07FBE138D903501A70235F6260885FA27028584A6D07FBE12",
         INIT_07 => x"7F01E702C6F17FFD04E703E702A7EF7FFD0000CC30E08E39D27FB7FF86016D84",
         INIT_08 => x"84A70520098D042420810D20608D0427F27F7D30E08E16345986028D1B86F27F",
         INIT_09 => x"270C81890027100D81382716817C0027101A815A271B81342708819635AF0017",
         INIT_0a => x"EF7FB66D205A34275DEF7FFC8F0016792619C15CEF7FFC45260A810F270B8124",
         INIT_0b => x"816E27598114273DC1F27FF656200000CC5820212750814CEF7FB662204A2C27",
         INIT_0c => x"224F812080F27F7F39F17FB70426F17F7D39F27F7F39F27FB704263D81312754",
         INIT_0d => x"508102A74C84E720C6EF7FB6168D0000CC1B20E12218C120C0F17F7FF17FF6ED",
         INIT_0e => x"EA2619C15C4FF02650814CEF7FFC3903E702A7EF7FFDF07FF64F39F27F7FF726",
         INIT_0f => x"7FF6F42650C15C84A702E7EF7FF72086EF7FF604E75F012519C15C04E6E78D5A"
      )
      port map (
         clk     => clk,
         en      => en(2),
         we      => we,
         rst     => rst,
         addr    => addr(8 downto 0),
         di      => wdata,
         do      => xdata(2)
      );

   ROM03: RAMB4_S8
      generic map (
         INIT_00 => x"FB035CFB0267FB0139F27FF702E7EF7FF75FE4205F03E7F07FF7082719C15CF0",
         INIT_01 => x"4DAFFA5051FA4C8FF847E7F84546F9423BFB1946FB1830FB1524FB1051FB0472",
         INIT_02 => x"0A0DFFFFFFFF7EF991F891F891F891F87EF9C5F95472F958DBF853E0FB5292F8",
         INIT_03 => x"000A0D4B04202D202045335320524F4620362E31204755423930535953000000",
         INIT_04 => x"3D53552020043D43502020043D5053202004202D20043F54414857043E040000",
         INIT_05 => x"432020043D422020043D412020043D50442020043D58492020043D5949202004",
         INIT_06 => x"C07F9F6E38F916D27FF7535FC07FCE103904315343565A4E4948464504203A43",
         INIT_07 => x"FF8CCC7FBE49584F4AAF80E64AAE431FCA7F9F6EC87F9F6EC67F9F6EC47F9F6E",
         INIT_08 => x"000000000000C27F9F6E42EE1F37F16E44AEC4EC10340822CE7FBC8B300F27FF",
         INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0a => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0b => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0c => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0d => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0e => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0f => x"D0FEDCFEECFEE8FEE4FEE0FEF0FEDCFE00000000000000000000000000000000"
      )
      port map (
         clk     => clk,
         en      => en(3),
         we      => we,
         rst     => rst,
         addr    => addr(8 downto 0),
         di      => wdata,
         do      => xdata(3)
      );

   rom_glue: process (cs, rw, addr, xdata)
   begin
      en <= (others=>'0');
      case addr(10 downto 9) is
      when "00" =>
         en(0)  <= cs;
         rdata  <= xdata(0);
      when "01" =>
         en(1)  <= cs;
         rdata  <= xdata(1);
      when "10" =>
         en(2)  <= cs;
         rdata  <= xdata(2);
      when "11" =>
         en(3)  <= cs;
         rdata  <= xdata(3);
      when others =>
         null;
      end case;
      we <= not rw;
   end process;
end architecture rtl;

