--=========================================================================
--
--  S Y N T H E Z I A B L E    SBUG - Monitor ROM for System09.
--
--=========================================================================
--
--  www.OpenCores.Org - September 2003
--  This core adheres to the GNU public license  
-- 
--         FILE NAME: sbug_rom2k_slice.vhd
--       ENTITY NAME: mon_rom
-- ARCHITECTURE NAME: rtl
--           VERSION: 1.0
--            AUTHOR: John E. Kent
--              DATE: 15 December 2002
--      DEPENDENCIES: ieee.Std_Logic_1164
--                    ieee.std_logic_unsigned
--                    ieee.std_logic_arith
--       DESCRIPTION: 2048 byte x 8 bit ROM Monitor program
--                    for the System09 using distributed RAM.
--                    ROM  sits at $F800
--                    ACIA sits at $E004
--                    DAT  sits at $FFF0
--         REVISIONS: 28th Jan 2007 
--                    Made entity compatible with Block RAM version
--

library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_arith.all;
	use ieee.std_logic_unsigned.all;

library unisim;
	use unisim.vcomponents.all;

entity mon_rom is
    Port (
       clk   : in  std_logic;
       rst   : in  std_logic;
       cs    : in  std_logic;
       rw    : in  std_logic;
       addr  : in  std_logic_vector (10 downto 0);
       wdata : in  std_logic_vector (7 downto 0);
       rdata : out std_logic_vector (7 downto 0)
    );
end mon_rom;

architecture rtl of mon_rom is


  constant width   : integer := 8;

  constant memsize : integer := 2048;


  type rom_array is array(0 to memsize-1) of std_logic_vector(width-1 downto 0);



  constant rom_data : rom_array :=
(

"11111000",
"00010100",
"11111000",
"01100001",
"11111101",
"11001111",
"11111101",
"11001001",
"11111101",
"11011111",
"11111101",
"11101110",
"11111101",
"10111101",
"11111101",
"10110001",
"11111101",
"10101101",
"11111011",
"10000001",
"10001110",
"11111110",
"01001111",
"00010000",
"10001110",
"11011111",
"11000000",
"11000110",
"00010000",
"10100110",
"10000000",
"10100111",
"10100000",
"01011010",
"00100110",
"11111001",
"10001110",
"11100000",
"00000100",
"10111111",
"11011111",
"11100000",
"00010111",
"00000010",
"01111010",
"11000110",
"00001100",
"01101111",
"11100010",
"01011010",
"00100110",
"11111011",
"00110000",
"10001100",
"11011101",
"10101111",
"01101010",
"10000110",
"11010000",
"10100111",
"11100100",
"00011111",
"01000011",
"00010111",
"00000101",
"10111110",
"10001110",
"11111110",
"01011111",
"00010111",
"00000101",
"01110101",
"10001110",
"11011111",
"11010000",
"01001111",
"11000110",
"00001101",
"01101101",
"10000101",
"00100111",
"00000011",
"10001011",
"00000100",
"00011001",
"01011010",
"00101010",
"11110110",
"00010111",
"00000101",
"00100110",
"10001110",
"11111110",
"01110100",
"00010111",
"00000101",
"01011100",
"10001110",
"11111110",
"01111011",
"00010111",
"00000101",
"01000110",
"00010111",
"00000101",
"01100101",
"10000100",
"01111111",
"10000001",
"00001101",
"00100111",
"11110001",
"00011111",
"10001001",
"10000001",
"00100000",
"00101100",
"00001001",
"10000110",
"01011110",
"00010111",
"00000101",
"01110011",
"00011111",
"10011000",
"10001011",
"01000000",
"00010111",
"00000101",
"01101100",
"00010111",
"00000101",
"01100111",
"11000001",
"01100000",
"00101111",
"00000010",
"11000000",
"00100000",
"10001110",
"11111110",
"00010011",
"11100001",
"10000000",
"00100111",
"00001111",
"00110000",
"00000010",
"10001100",
"11111110",
"01001111",
"00100110",
"11110101",
"10001110",
"11111110",
"01111101",
"00010111",
"00000101",
"00011110",
"00100000",
"11000000",
"10101101",
"10010100",
"00100000",
"10111100",
"00011111",
"00110100",
"00111011",
"10001110",
"11111110",
"10000011",
"00010111",
"00000100",
"11111111",
"00010111",
"00000100",
"00010001",
"00010111",
"00000100",
"00011001",
"00010111",
"00000100",
"00100001",
"00010111",
"00000100",
"00101001",
"00010111",
"00000100",
"00110001",
"10001110",
"11111110",
"10000011",
"00010111",
"00000100",
"11101010",
"00010111",
"00000100",
"00110011",
"00010111",
"00000100",
"00111010",
"00010111",
"00000100",
"01000001",
"00010110",
"00000100",
"01001000",
"00010111",
"00000100",
"00100111",
"00010111",
"00000101",
"00010111",
"00010111",
"00000100",
"01010111",
"00101001",
"00000010",
"10101111",
"01001010",
"00111001",
"00010111",
"00000011",
"11101101",
"00010111",
"00000101",
"00001001",
"00010111",
"00000100",
"01001001",
"00101001",
"00000010",
"10101111",
"01001000",
"00111001",
"00010111",
"00000100",
"00000000",
"00010111",
"00000100",
"11111011",
"00010111",
"00000100",
"00111011",
"00101001",
"00000010",
"10101111",
"01000110",
"00111001",
"00010111",
"00000011",
"11100111",
"00010111",
"00000100",
"11101101",
"00010111",
"00000100",
"00101101",
"00101001",
"00000010",
"10101111",
"01000100",
"00111001",
"00010111",
"00000011",
"11001110",
"00010111",
"00000100",
"11011111",
"00010111",
"00000100",
"00110000",
"00101001",
"00000010",
"10100111",
"01000011",
"00111001",
"00010111",
"00000011",
"11110101",
"00010111",
"00000100",
"11010001",
"00010111",
"00000100",
"00100010",
"00101001",
"00000010",
"10100111",
"01000010",
"00111001",
"00010111",
"00000011",
"11011101",
"00010111",
"00000100",
"11000011",
"00010111",
"00000100",
"00010100",
"00101001",
"00000010",
"10100111",
"01000001",
"00111001",
"00010111",
"00000011",
"11100011",
"00010111",
"00000100",
"10110101",
"00010111",
"00000100",
"00000110",
"00101001",
"00000100",
"10001010",
"10000000",
"10100111",
"11000100",
"00111001",
"00010111",
"00000011",
"11101011",
"00101001",
"00101101",
"00011111",
"00010010",
"10001110",
"11111110",
"10000011",
"00010111",
"00000100",
"01011111",
"00011111",
"00100001",
"00010111",
"00000100",
"00100110",
"00010111",
"00000100",
"10010110",
"10100110",
"10100100",
"00010111",
"00000100",
"00100110",
"00010111",
"00000100",
"10001110",
"00010111",
"00000011",
"11011111",
"00101000",
"00010001",
"10000001",
"00001000",
"00100111",
"11100001",
"10000001",
"00011000",
"00100111",
"11011101",
"10000001",
"01011110",
"00100111",
"00010111",
"10000001",
"00001101",
"00100110",
"00001111",
"00111001",
"10100111",
"10100100",
"10100001",
"10100100",
"00100111",
"00001000",
"00010111",
"00000100",
"01101111",
"10000110",
"00111111",
"00010111",
"00000100",
"01101100",
"00110001",
"00100001",
"00100000",
"11000010",
"00110001",
"00111111",
"00100000",
"10111110",
"00010111",
"00000011",
"00110101",
"00011111",
"00110010",
"10001110",
"11011111",
"11000000",
"00110000",
"00011111",
"00100000",
"00000101",
"00010111",
"00000011",
"10001011",
"00101001",
"00000110",
"00110100",
"00100000",
"10101100",
"11100001",
"00100100",
"00000001",
"00111001",
"00011111",
"00010000",
"11000011",
"00000000",
"00010000",
"11000100",
"11110000",
"00110100",
"00000110",
"00011111",
"00100000",
"11000100",
"11110000",
"00011111",
"00000001",
"10101100",
"11100100",
"00100111",
"00000101",
"00010111",
"00000100",
"00100111",
"00100111",
"00000011",
"00110010",
"01100010",
"00111001",
"00110100",
"00010000",
"10001110",
"11111110",
"10000011",
"00010111",
"00000011",
"11101000",
"10101110",
"11100100",
"00010111",
"00000011",
"10101111",
"11000110",
"00010000",
"10100110",
"10000000",
"00010111",
"00000011",
"10110000",
"00010111",
"00000100",
"00011000",
"01011010",
"00100110",
"11110101",
"00010111",
"00000100",
"00010000",
"10101110",
"11100001",
"11000110",
"00010000",
"10100110",
"10000000",
"10000001",
"00100000",
"00100101",
"00000100",
"10000001",
"01111110",
"00100011",
"00000010",
"10000110",
"00101110",
"00010111",
"00000100",
"00000001",
"01011010",
"00100110",
"11101110",
"00100000",
"10111111",
"01101111",
"11100010",
"01101111",
"11100010",
"00010111",
"00000011",
"00101011",
"00110100",
"00110000",
"00101001",
"01111011",
"10101100",
"01100010",
"00100101",
"01110111",
"00010111",
"00000011",
"11101000",
"00011111",
"00100000",
"11100011",
"01100100",
"00110100",
"00000100",
"10101011",
"11100000",
"10100111",
"10100000",
"00010000",
"10101100",
"11100100",
"00100101",
"11110001",
"00010000",
"10101110",
"01100010",
"00011111",
"00100000",
"11100011",
"01100100",
"00110100",
"00000010",
"11101011",
"11100000",
"11101000",
"10100000",
"00100111",
"00111100",
"10001110",
"11111110",
"10000011",
"00010111",
"00000011",
"10000101",
"00110000",
"00111111",
"00010111",
"00000011",
"01001100",
"00110100",
"00010000",
"10001110",
"11111110",
"10100001",
"00010111",
"00000011",
"10001000",
"00110101",
"00010000",
"00010111",
"00000001",
"01000111",
"00010111",
"00000011",
"01010000",
"00010111",
"00000011",
"00111001",
"10001110",
"11111110",
"10000111",
"00010111",
"00000011",
"01110111",
"10101110",
"01100100",
"00010111",
"00000011",
"00101110",
"10001110",
"11111110",
"10001111",
"00010111",
"00000011",
"01101100",
"00011111",
"10011000",
"10001110",
"11111110",
"10100110",
"00010111",
"00000011",
"00111110",
"00010111",
"00000011",
"10000011",
"00100110",
"00011010",
"00010000",
"10101100",
"11100100",
"00100101",
"10110011",
"10000110",
"00101011",
"00010111",
"00000011",
"10000110",
"00010111",
"00000011",
"01110100",
"00100110",
"00001011",
"00010000",
"10101110",
"01100010",
"01101100",
"01100101",
"00100110",
"10010000",
"01101100",
"01100100",
"00100110",
"10001100",
"00110010",
"01100110",
"00111001",
"00010111",
"00000010",
"10110001",
"00101001",
"00011110",
"10001100",
"11011111",
"11000000",
"00100100",
"00011010",
"00110100",
"00010000",
"10001110",
"11111111",
"11111111",
"10001101",
"01010101",
"00110101",
"00010000",
"00100111",
"00001111",
"10100110",
"10000100",
"10000001",
"00111111",
"00100111",
"00001001",
"10100111",
"10100000",
"10101111",
"10100100",
"10000110",
"00111111",
"10100111",
"10000100",
"00111001",
"00010111",
"00000011",
"01001010",
"10000110",
"00111111",
"00010110",
"00000011",
"01000111",
"00010000",
"10001110",
"11011111",
"11100011",
"11000110",
"00001000",
"10001101",
"00011000",
"01011010",
"00100110",
"11111011",
"00111001",
"00011111",
"01000011",
"10101110",
"01001010",
"00110000",
"00011111",
"10001101",
"00100110",
"00100111",
"00000100",
"10101111",
"01001010",
"10001101",
"00000110",
"00010111",
"11111101",
"11100100",
"00010110",
"11111101",
"10011010",
"10101110",
"00100001",
"10001100",
"11011111",
"11000000",
"00100100",
"00001010",
"10100110",
"10000100",
"10000001",
"00111111",
"00100110",
"00000100",
"10100110",
"10100100",
"10100111",
"10000100",
"10000110",
"11111111",
"10100111",
"10100000",
"10100111",
"10100000",
"10100111",
"10100000",
"00111001",
"00010000",
"10001110",
"11011111",
"11100011",
"11000110",
"00001000",
"10100110",
"10100000",
"10101100",
"10100001",
"00100111",
"00000100",
"01011010",
"00100110",
"11110111",
"00111001",
"00110001",
"00111101",
"00111001",
"10000110",
"11011110",
"10110111",
"11110000",
"00100100",
"10000110",
"11111111",
"10110111",
"11110000",
"00010100",
"10110111",
"11110000",
"00010000",
"10110111",
"11110000",
"00010101",
"10110111",
"11110000",
"00010110",
"01111101",
"11110000",
"00010000",
"10000110",
"11011000",
"10110111",
"11110000",
"00100000",
"00010111",
"00000000",
"10010111",
"10110110",
"11110000",
"00100000",
"00101011",
"11111011",
"10000110",
"00001001",
"10110111",
"11110000",
"00100000",
"00010111",
"00000000",
"10001010",
"10110110",
"11110000",
"00100000",
"10000101",
"00000001",
"00100110",
"11111001",
"10000101",
"00010000",
"00100110",
"11001010",
"10001110",
"11000000",
"00000000",
"10001101",
"01010010",
"10001010",
"00010000",
"10110111",
"11110000",
"01000000",
"00011111",
"00010000",
"01000011",
"01010011",
"11111101",
"11110000",
"00000000",
"10001110",
"11111110",
"11111111",
"10111111",
"11110000",
"00000010",
"10000110",
"11111111",
"10110111",
"11110000",
"00010000",
"10000110",
"11111110",
"10110111",
"11110000",
"00010100",
"10000110",
"00000001",
"10110111",
"11110000",
"00100010",
"10000110",
"10001100",
"10110111",
"11110000",
"00100000",
"10001101",
"01010010",
"01011111",
"00110100",
"00000100",
"01011111",
"01111101",
"11110000",
"00010000",
"00101010",
"00001010",
"01011010",
"00100110",
"11111000",
"00110101",
"00000100",
"01011010",
"00100110",
"11110000",
"00100000",
"10001010",
"00110101",
"00000100",
"10110110",
"11110000",
"00100000",
"10000101",
"00011100",
"00100111",
"00000001",
"00111001",
"11000110",
"11011110",
"11110111",
"11110000",
"00100100",
"10001110",
"11000000",
"00000000",
"10101111",
"01001010",
"00011111",
"00110100",
"00111011",
"00110100",
"00110110",
"10100110",
"01100010",
"01000100",
"01000100",
"01000100",
"01000100",
"00010000",
"10001110",
"11011111",
"11010000",
"11100110",
"10100110",
"01010100",
"01010100",
"01010100",
"01010100",
"11100111",
"11100100",
"11100110",
"10100110",
"01010011",
"01011000",
"01011000",
"01011000",
"01011000",
"10100110",
"01100010",
"10000100",
"00001111",
"10100111",
"01100010",
"11101010",
"01100010",
"11100111",
"01100010",
"00110101",
"00110110",
"00111001",
"00110100",
"00000100",
"11000110",
"00100000",
"01011010",
"00100110",
"11111101",
"00110101",
"00000100",
"00111001",
"01111101",
"11100000",
"00011000",
"01111111",
"11100000",
"00010100",
"11000110",
"00000011",
"10001110",
"00000000",
"00000000",
"00110000",
"00000001",
"10001100",
"00000000",
"00000000",
"00100110",
"11111001",
"01011010",
"00100110",
"11110110",
"10000110",
"00001111",
"10110111",
"11100000",
"00011000",
"10001101",
"00110111",
"11110110",
"11100000",
"00011000",
"11000101",
"00000001",
"00100110",
"11111001",
"10000110",
"00000001",
"10110111",
"11100000",
"00011010",
"10001101",
"00101001",
"10000110",
"10001100",
"10110111",
"11100000",
"00011000",
"10001101",
"00100010",
"10001110",
"11000000",
"00000000",
"00100000",
"00001001",
"11000101",
"00000010",
"00100111",
"00000101",
"10110110",
"11100000",
"00011011",
"10100111",
"10000000",
"11110110",
"11100000",
"00011000",
"11000101",
"00000001",
"00100110",
"11110000",
"11000101",
"00101100",
"00100111",
"00000001",
"00111001",
"10001110",
"11000000",
"00000000",
"10101111",
"01001010",
"00011111",
"00110100",
"00111011",
"11000110",
"00100000",
"01011010",
"00100110",
"11111101",
"00111001",
"10000110",
"00010001",
"00010111",
"00000001",
"11011101",
"01111111",
"11011111",
"11100010",
"00010111",
"00000001",
"10101101",
"10000001",
"01010011",
"00100110",
"11111001",
"00010111",
"00000001",
"10100110",
"10000001",
"00111001",
"00100111",
"00111101",
"10000001",
"00110001",
"00100110",
"11110001",
"00010111",
"00000001",
"00010111",
"00110100",
"00000010",
"00101001",
"00100110",
"00010111",
"00000000",
"11111111",
"00101001",
"00100001",
"00110100",
"00010000",
"11100110",
"11100000",
"11101011",
"11100000",
"11101011",
"11100100",
"01101010",
"11100100",
"01101010",
"11100100",
"00110100",
"00000100",
"00010111",
"00000000",
"11111101",
"00110101",
"00000100",
"00101001",
"00001100",
"00110100",
"00000010",
"11101011",
"11100000",
"01101010",
"11100100",
"00100111",
"00000101",
"10100111",
"10000000",
"00100000",
"11101011",
"01011111",
"00110101",
"00000010",
"11000001",
"11111111",
"00100111",
"10110010",
"10000110",
"00111111",
"00010111",
"00000001",
"10001111",
"01110011",
"11011111",
"11100010",
"10000110",
"00010011",
"00010110",
"00000001",
"10000111",
"01101111",
"11100010",
"00010111",
"00000000",
"10111000",
"00110100",
"00110000",
"00101001",
"01001010",
"10101100",
"01100010",
"00100101",
"01000110",
"00110000",
"00000001",
"10101111",
"11100100",
"10000110",
"00010010",
"00010111",
"00000001",
"01110001",
"11101100",
"11100100",
"10100011",
"01100010",
"00100111",
"00000110",
"00010000",
"10000011",
"00000000",
"00100000",
"00100011",
"00000010",
"11000110",
"00100000",
"11100111",
"01100100",
"10001110",
"11111110",
"11101011",
"00010111",
"00000001",
"00011010",
"11001011",
"00000011",
"00011111",
"10011000",
"00010111",
"00000000",
"11100111",
"10101110",
"01100010",
"00010111",
"00000000",
"11011010",
"11101011",
"01100010",
"11101011",
"01100011",
"11101011",
"10000100",
"10100110",
"10000000",
"00010111",
"00000000",
"11010111",
"01101010",
"01100100",
"00100110",
"11110101",
"01010011",
"00011111",
"10011000",
"00010111",
"00000000",
"11001101",
"10101111",
"01100010",
"10101100",
"11100100",
"00100110",
"11000011",
"10000110",
"00010100",
"00010111",
"00000001",
"00101111",
"00110010",
"01100101",
"00111001",
"10001110",
"11111110",
"10101110",
"00010111",
"00000000",
"11110101",
"00011111",
"00110001",
"00010110",
"00000000",
"10101100",
"10001110",
"11111110",
"10111010",
"00010111",
"00000000",
"11101010",
"10101110",
"01001000",
"00010110",
"00000000",
"10100001",
"10001110",
"11111110",
"11001100",
"00010111",
"00000000",
"11011111",
"10100110",
"01000011",
"00010110",
"00000000",
"10011110",
"10001110",
"11111110",
"11000110",
"00010111",
"00000000",
"11010100",
"10101110",
"01000100",
"00010110",
"00000000",
"10001011",
"10001110",
"11111110",
"11000000",
"00010111",
"00000000",
"11001001",
"10101110",
"01000110",
"00010110",
"00000000",
"10000000",
"10001110",
"11111110",
"10110100",
"00010111",
"00000000",
"10111110",
"10101110",
"01001010",
"00100000",
"01110110",
"10001110",
"11111110",
"11010010",
"00010111",
"00000000",
"10110100",
"10100110",
"01000001",
"00100000",
"01110100",
"10001110",
"11111110",
"11010111",
"00010111",
"00000000",
"10101010",
"10100110",
"01000010",
"00100000",
"01101010",
"10001110",
"11111110",
"11011100",
"00010111",
"00000000",
"10100000",
"10100110",
"11000100",
"10001110",
"11111110",
"11100011",
"00100000",
"01110011",
"10001101",
"00001001",
"00101001",
"01001110",
"00011111",
"00010010",
"10000110",
"00101101",
"00010111",
"00000000",
"10111111",
"10001101",
"00001111",
"00101001",
"01000011",
"00011111",
"00000001",
"10001101",
"00001001",
"00101001",
"00111101",
"00110100",
"00010000",
"10100111",
"01100001",
"00110101",
"00010000",
"00111001",
"10001101",
"00010001",
"00101001",
"00110010",
"01001000",
"01001000",
"01001000",
"01001000",
"00011111",
"10001001",
"10001101",
"00000111",
"00101001",
"00101000",
"00110100",
"00000100",
"10101011",
"11100000",
"00111001",
"10001101",
"01101111",
"10000001",
"00110000",
"00100101",
"00011101",
"10000001",
"00111001",
"00100010",
"00000011",
"10000000",
"00110000",
"00111001",
"10000001",
"01000001",
"00100101",
"00010010",
"10000001",
"01000110",
"00100010",
"00000011",
"10000000",
"00110111",
"00111001",
"10000001",
"01100001",
"00100101",
"00000111",
"10000001",
"01100110",
"00100010",
"00000011",
"10000000",
"01010111",
"00111001",
"00011010",
"00000010",
"00111001",
"00110100",
"00010000",
"00110101",
"00000010",
"10001101",
"00000010",
"00110101",
"00000010",
"00110100",
"00000010",
"01000100",
"01000100",
"01000100",
"01000100",
"10001101",
"00000100",
"00110101",
"00000010",
"10000100",
"00001111",
"10001011",
"00110000",
"10000001",
"00111001",
"00101111",
"00000010",
"10001011",
"00000111",
"00100000",
"01010111",
"00110100",
"00000010",
"11000110",
"00001000",
"10100110",
"10000000",
"01101000",
"11100100",
"00100101",
"00000010",
"10000110",
"00101101",
"10001101",
"01001001",
"10001101",
"01000101",
"01011010",
"00100110",
"11110001",
"00110101",
"00000010",
"00111001",
"10001101",
"00000010",
"00100000",
"00001100",
"00110100",
"00010000",
"10001110",
"11111110",
"01110101",
"10001101",
"00000101",
"00110101",
"00010000",
"00111001",
"10001101",
"00110001",
"10100110",
"10000000",
"10000001",
"00000100",
"00100110",
"11111000",
"00111001",
"01111101",
"11011111",
"11100010",
"00100111",
"00000110",
"10001101",
"00000100",
"10000100",
"01111111",
"00100000",
"00011111",
"00110100",
"00010000",
"10111110",
"11011111",
"11100000",
"10100110",
"10000100",
"10000101",
"00000001",
"00100111",
"11111010",
"10100110",
"00000001",
"00110101",
"00010000",
"00111001",
"00110100",
"00000010",
"10100110",
"10011111",
"11011111",
"11100000",
"10000101",
"00000001",
"00110101",
"00000010",
"00111001",
"10001101",
"00000000",
"10000110",
"00100000",
"00110100",
"00010010",
"10111110",
"11011111",
"11100000",
"10100110",
"10000100",
"10000101",
"00000010",
"00100111",
"11111010",
"00110101",
"00000010",
"10100111",
"00000001",
"00110101",
"00010000",
"00111001",
"10111110",
"11011111",
"11100000",
"10000110",
"00000011",
"10100111",
"10000100",
"10000110",
"00010001",
"10100111",
"10000100",
"01101101",
"00000001",
"10000110",
"11111111",
"10110111",
"11011111",
"11100010",
"00111001",
"00000001",
"11111001",
"00100011",
"00000010",
"11111001",
"00010101",
"00000011",
"11111001",
"00110001",
"00000100",
"11111001",
"00000111",
"00010000",
"11111000",
"11001111",
"00010101",
"11111000",
"11011101",
"00011000",
"11111000",
"11111001",
"00011001",
"11111000",
"11101011",
"01000010",
"11111010",
"01111011",
"01000100",
"11111010",
"11110100",
"01000101",
"11111001",
"10010110",
"01000111",
"11111000",
"10100101",
"01001100",
"11111100",
"00001100",
"01001101",
"11111001",
"01000001",
"01010000",
"11111100",
"01100111",
"01010001",
"11111001",
"11110010",
"01010010",
"11111000",
"10101000",
"01010011",
"11111001",
"10001010",
"01010101",
"11111011",
"10110011",
"01011000",
"11111010",
"10100111",
"11111010",
"10110011",
"11111000",
"10100111",
"11111000",
"10100111",
"11111000",
"10100111",
"11111000",
"10100111",
"11111010",
"10110011",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"00001101",
"00001010",
"00000000",
"00000000",
"00000000",
"01010011",
"00101101",
"01000010",
"01010101",
"01000111",
"00100000",
"00110001",
"00101110",
"00111000",
"00100000",
"00101101",
"00100000",
"00000100",
"01001011",
"00001101",
"00001010",
"00000000",
"00000000",
"00000000",
"00000100",
"00111110",
"00000100",
"01010111",
"01001000",
"01000001",
"01010100",
"00111111",
"00000100",
"00100000",
"00101101",
"00100000",
"00000100",
"00101100",
"00100000",
"01010000",
"01000001",
"01010011",
"01010011",
"00100000",
"00000100",
"00101100",
"00100000",
"01000010",
"01001001",
"01010100",
"01010011",
"00100000",
"01001001",
"01001110",
"00100000",
"01000101",
"01010010",
"01010010",
"01001111",
"01010010",
"00111010",
"00100000",
"00000100",
"00100000",
"00111101",
"00111110",
"00100000",
"00000100",
"00110111",
"00110110",
"00110101",
"00110100",
"00110011",
"00110010",
"00110001",
"00110000",
"00100000",
"00100000",
"01010011",
"01010000",
"00111101",
"00000100",
"00100000",
"00100000",
"01010000",
"01000011",
"00111101",
"00000100",
"00100000",
"00100000",
"01010101",
"01010011",
"00111101",
"00000100",
"00100000",
"00100000",
"01001001",
"01011001",
"00111101",
"00000100",
"00100000",
"00100000",
"01001001",
"01011000",
"00111101",
"00000100",
"00100000",
"00100000",
"01000100",
"01010000",
"00111101",
"00000100",
"00100000",
"00100000",
"01000001",
"00111101",
"00000100",
"00100000",
"00100000",
"01000010",
"00111101",
"00000100",
"00100000",
"00100000",
"01000011",
"01000011",
"00111010",
"00100000",
"00000100",
"01000101",
"01000110",
"01001000",
"01001001",
"01001110",
"01011010",
"01010110",
"01000011",
"01010011",
"00110001",
"00000100",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"00000000",
"00000000",
"00000000",
"10001110",
"11111111",
"11110000",
"10000110",
"00001111",
"10100111",
"10000000",
"01001010",
"00100110",
"11111011",
"10000110",
"11110000",
"10100111",
"10000100",
"10001110",
"11010000",
"10100000",
"00010000",
"10001110",
"01010101",
"10101010",
"11101110",
"10000100",
"00010000",
"10101111",
"10000100",
"00010000",
"10101100",
"10000100",
"00100111",
"00001011",
"00110000",
"10001001",
"11110000",
"00000000",
"10001100",
"11110000",
"10100000",
"00100110",
"11101101",
"00100000",
"11010110",
"11101111",
"10000100",
"00011111",
"00010000",
"01000011",
"01000100",
"01000100",
"01000100",
"01000100",
"10110111",
"11111111",
"11111101",
"00010000",
"11001110",
"11011111",
"11000000",
"00010000",
"10001110",
"11011111",
"11010000",
"10100111",
"00101101",
"01101111",
"00101110",
"10000110",
"11110000",
"10100111",
"00101111",
"10000110",
"00001100",
"01101111",
"10100110",
"01001010",
"00101010",
"11111011",
"00110000",
"10001001",
"11110000",
"00000000",
"10001100",
"11110000",
"10100000",
"00100111",
"00100010",
"11101110",
"10000100",
"00010000",
"10001110",
"01010101",
"10101010",
"00010000",
"10101111",
"10000100",
"00010000",
"10101100",
"10000100",
"00100110",
"11101001",
"11101111",
"10000100",
"00010000",
"10001110",
"11011111",
"11010000",
"00011111",
"00010000",
"01000100",
"01000100",
"01000100",
"01000100",
"00011111",
"10001001",
"10001000",
"00001111",
"10100111",
"10100101",
"00100000",
"11010101",
"10000110",
"11110001",
"00010000",
"10001110",
"11011111",
"11010000",
"10100111",
"00101110",
"10000110",
"00001100",
"11100110",
"10100110",
"00100110",
"00000101",
"01001010",
"00101010",
"11111001",
"00100000",
"00010100",
"01101111",
"10100110",
"11100111",
"00101100",
"01001111",
"00011111",
"00100001",
"11100110",
"10100110",
"00100111",
"00000100",
"01101111",
"10100110",
"11100111",
"10000000",
"01001100",
"10000001",
"00001100",
"00101101",
"11110011",
"10001110",
"11111111",
"11110000",
"11000110",
"00010000",
"10100110",
"10100000",
"10100111",
"10000000",
"01011010",
"00100110",
"11111001",
"01010011",
"11110111",
"11011111",
"11100010",
"00010110",
"11111000",
"01100010",
"01101110",
"10011111",
"11011111",
"11000000",
"01101110",
"10011111",
"11011111",
"11000100",
"01101110",
"10011111",
"11011111",
"11000110",
"01101110",
"10011111",
"11011111",
"11001000",
"01101110",
"10011111",
"11011111",
"11001010",
"00011111",
"01000011",
"10101110",
"01001010",
"11100110",
"10000000",
"10101111",
"01001010",
"01001111",
"01011000",
"01001001",
"10111110",
"11011111",
"11001100",
"10001100",
"11111111",
"11111111",
"00100111",
"00001111",
"00110000",
"10001011",
"10111100",
"11011111",
"11001110",
"00100010",
"00001000",
"00110100",
"00010000",
"11101100",
"11000100",
"10101110",
"01000100",
"01101110",
"11110001",
"00110111",
"00011111",
"11101110",
"01000010",
"01101110",
"10011111",
"11011111",
"11000010",
"11111111",
"10110010",
"11111111",
"11000110",
"11111111",
"10110110",
"11111111",
"10111010",
"11111111",
"10111110",
"11111111",
"11000010",
"11111111",
"10110010",
"11111111",
"00000000"
);
begin

   rdata <= rom_data(conv_integer(addr)); 


end architecture;

