    INIT_00 => x"54C74AD354C7B7D201BCC2B4C6FEF77BC2D4C85BBCC289C6AEC9E6C77EE2D6C5",
    INIT_01 => x"5D45534C45057DD554C7FAF76EC2AFC046C736F898C273D35D4E454854057DD5",
    INIT_02 => x"46C768F898C273D35D4649037DD554C7FAF76EC2AFC0C9C746C750F898C273D3",
    INIT_03 => x"F7FAF76EC2AEC9E6C77BF898C273D35D4441454841067DD5FAF76EC2AEC9E6C7",
    INIT_04 => x"C0BD5D44414548415B0701EEF57EC0F7F700BCC2FFC0BD5D45534C455B0601DA",
    INIT_05 => x"C2FFC0BD534D020202F17EC089F892C0FFC0BD5D46495B040185F07EC089F8FF",
    INIT_06 => x"0188A8F813D17EC0C6F83DC3D0F83DC3D4F807C300BCC212BCC2D8F825C300BC",
    INIT_07 => x"B4C6D9D3D6C500BCC2FFC0BD4745520309BCF77EC03300CBC200BCC2FFC0BD23",
    INIT_08 => x"F8E6D4E8E342D5DBC707F93DC3DDC643C9D1C600C8FBD6B4C617F925C300BCC2",
    INIT_09 => x"BD2950440308C5F67EC0E1F8FF00AFC2FFC0BD4745524C4C4106084AF77EC0E1",
    INIT_0a => x"73F77EC0D0D68900AFC200C8FFC0BD2923020882F87EC03300CBC210BCC2FFC0",
    INIT_0b => x"18C4FFC0BD5D5B02084EF97EC08D00AFC23300CBC220BCC2FFC0BD2943500308",
    INIT_0c => x"7EC0D7C910BCC2B8D6D4C88000AFC237C99D00AFC2E6C7A0F97BC2D4C820BCC2",
    INIT_0d => x"C4FDCC00BCC2FDCCFFC0BD4649028896F886EB7EC09F00AFC23300CBC220BCC2",
    INIT_0e => x"F4CDEB7EC0B5F920BCC2FFC0BD44414548410588B2F9A4EB7EC0BFCD06BCC2A7",
    INIT_0f => x"C8B8D6ABC886D6E6C7E0C9F2C7A7C495D406BCC2D3CDFFC0BD4E4548540488E5",
    INIT_10 => x"04EC7EC0BFCD07BCC2A7C4FFC0BD4E4947454205883BF9EBEB7EC01DC6B9C900",
    INIT_11 => x"D6E6C7E0C9AEC9A7C4FDCC00C895D407BCC2D3CDFFC0BD4C49544E55058878F9",
    INIT_12 => x"3EEC7EC029FA20BCC2FFC0BD4E49414741058823FA23EC7EC0FDCCB8D6ABC886",
    INIT_13 => x"45504552068841F654EC7EC0E7F912CE01BCC2D3F9FFC0BD45534C4504885AF3",
    INIT_14 => x"12CE01BCC2B5F9FFC0BD454C49485705884EFAB8EB7EC0E7F954FAFFC0BD5441",
    INIT_15 => x"2D444345530B0690FA7EC0ACDA7BF99CE044E0FFC0BD5458454E0408D0F77EC0",
    INIT_16 => x"484749482D535345524444412D44434553110626F940B152C1BD535554415453",
    INIT_17 => x"530A06B9F800B252C1BD455341422D4D41522D444345530D06CDF941B152C1BD",
    INIT_18 => x"544154532D444345532E0C06E2F97EC002D2A7C4FFC0BD54524154532D444345",
    INIT_19 => x"088DD5B5F9ABC837C901BCC2E6C789C6C6FA203A44434553068DD5FFC0BD5355",
    INIT_1a => x"C903BCC288C901BCC2E7F920444550504F5453088DD568FA20474E494E4E5552",
    INIT_1b => x"D5B5F9D4C801BCC2E6C7E7F9474E494E4E5552078DD5B5F9D4C800BCC2E6C737",
    INIT_1c => x"F9D4C803BCC2E7F94347028DD5B5F9D4C802BCC2E6C7E7F94445544C4148068D",
    INIT_1d => x"BD454741502D444345532E0A0610F27EC059CFE7F94E574F4E4B4E55078DD5B5",
    INIT_1e => x"4553080659F17EC02CC6CCC406F50001AFC2F6FA77D295C6CCC41DC6E0FAFFC0",
    INIT_1f => x"6E61206874726F467369614D0F000000007EC002D2A7C4FFC0BD444E452D4443",
    INIT_20 => x"6B636174530F03FCFCFF776F6C667265766F206B636174530EEFFBFDFF313036",
    INIT_21 => x"6E4F0E2AFCF2FF646E69662074276E61430A16FCF3FF776F6C667265646E7520",
    INIT_22 => x"450C4CFCF0FF6465746365746F72500939FCF1FF676E696C69706D6F6320796C",
    INIT_23 => x"FF726F727265206572757463757274530F5AFCEAFF7475706E6920666F20646E",
    INIT_24 => x"6E2064696C61766E49157FFCE0FF747075727265746E6920726573550E6BFCE4",
    INIT_25 => x"766F20726564726F206863726165531592FCCFFF746E656D7567726120656D61",
    INIT_26 => x"6F6C667265646E7520726564726F2068637261655316ACFCCEFF776F6C667265",
    INIT_27 => x"72207369204553414218E1FCC2FF3F73696874207327746168570CC6FCC3FF77",
    INIT_28 => x"72646461206C6167656C6C4917F2FCC1FF6C616D69636564206F742074657365",
    INIT_29 => x"00000000000000000000000000000000E2C000000065646F6D20676E69737365",
    INIT_2a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2f => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3f => x"5EF1640061005E005B005800550000C000000000000000000000000000000000",
