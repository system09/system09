--
-- SYS09BUG Monitor Program
-- v1.0 - 21 November 2006 - John Knet
--
-- v1.1 - 22 december 2006 - John Kent
--        made into 4K ROM/RAM.
-- 
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
library unisim;
	use unisim.vcomponents.all;

entity mon_rom is
    Port (
       clk   : in  std_logic;
		 rst   : in  std_logic;
		 cs    : in  std_logic;
		 rw    : in  std_logic;
       addr  : in  std_logic_vector (11 downto 0);
       rdata : out std_logic_vector (7 downto 0);
       wdata : in  std_logic_vector (7 downto 0)
    );
end mon_rom;

architecture rtl of mon_rom is

  signal we     : std_logic;
  signal cs0    : std_logic;
  signal cs1    : std_logic;
  signal dp0    : std_logic;
  signal dp1    : std_logic;
  signal rdata0 : std_logic_vector(7 downto 0);
  signal rdata1 : std_logic_vector(7 downto 0);


begin

  ROM0 : RAMB16_S9
    generic map ( 
    INIT_00 => x"3FF13FF13FF141F119F152F052F052F03FF13FF13FF13FF13FF141F119F1BDF7",
    INIT_01 => x"7AF152F052F052F052F052F052F052F052F052F052F052F052F052F03FF13FF1",
    INIT_02 => x"6E34DE9F6E32DE9F6E39FE1C5D5F52F052F052F04EF24EF24EF24EF249F2E9F1",
    INIT_03 => x"0FC630350826FF8185A62ADE8E1EDEF703E6303438DE9F6E390127078D36DE9F",
    INIT_04 => x"6E3ADE9F6E3035F9265AA0A780A614C632DE8E108B3002F08E3D14C639011A5D",
    INIT_05 => x"6E39EA2604814C1EDEB640DE9FAD0425BC8D1BDE8E1EDEB74F3EDE9F6E3CDE9F",
    INIT_06 => x"F084C5AB1FDEB62EDECEC5E61EDEF62ADECE501A22DEB7A81F44DE9F6E42DE9F",
    INIT_07 => x"B70F88008639031F5F008B0F841FDEB6F0FFB7E0AB0F840F88018020DEB6E2A7",
    INIT_08 => x"FF17EAFF17703439011A5D40C639041AFE1C20DEF71FDEB7398A1F22DEB6F0FF",
    INIT_09 => x"5FF0355FF9265A80A7A0A65F46DE8E10CBFF17F9265AA0A7C0A65F46DE8E10A6",
    INIT_0a => x"80A65F46DE8E10BAFF16032700C1072701C1C5E61EDEF62ADECEC2FF17703439",
    INIT_0b => x"DE7F02340434F0355F84FF17F9265AC0A7A0A65F46DE8E105FFF17F9265AA0A7",
    INIT_0c => x"2485F2BD02353D2485F2BD0235442485F2BD1EDEB64C2485F2BD738622DE7F21",
    INIT_0d => x"F2BD02341B2467F2BDEB265A21DE7C032422DEB722DEBB80A7302467F2BD5F36",
    INIT_0e => x"85F2BD1586092010C60D205F032485F2BD06860E2621DEB3100235891F142467",
    INIT_0f => x"85F2BD1EDEB6DD2485F2BD728622DE7F21DE7F02340434395D21DEF709C6F524",
    INIT_10 => x"032422DEB722DEBBBF2485F2BD80A65FC72485F2BD0235CE2485F2BD0235D524",
    INIT_11 => x"5F032606819C2467F2BDA12485F2BD22DEB6A92485F2BD21DEB6EB265A21DE7C",
    INIT_12 => x"205F03260681072467F2BD0C2485F2BD5186395D21DEF6395D21DEF70AC60220",
    INIT_13 => x"B035EE261F30F6263F310A254700E0B6E2048E10E8038E3034395D011A10C604",
    INIT_14 => x"35ED261F30F5263F310C25474700E0B6E2048E10E8038E02343034B03501E0B6",
    INIT_15 => x"2E2E2E6B7369644D415220676E6974616D726F460D0AB03501E0B70235B03502",
    INIT_16 => x"AAF28E04202164657461636F6C6C6120746F6E206B7369646D6152040D0A0420",
    INIT_17 => x"BD1BDE8E1EDEF7396AF4BDC2F28EF52604C15C0C27018185A65F2ADE8E6AF4BD",
    INIT_18 => x"4C20DEB684A71FDEB646DE8E20DEB701861FDE7FFB265A80A75F4F46DE8E6CF0",
    INIT_19 => x"B70186D7260F8120DEB620DE7C5BF0BD20DEF61FDEB601A70186846C04260F81",
    INIT_1a => x"C6BF86016F846F46DE8E57F0BD0EC6BF8646DE8EC826C0811FDEB61FDE7C20DE",
    INIT_1b => x"03C64F46DE8E5BF0BD0EC64F016F846F46DE8E57F0BD0EC64F46DE8E5BF0BD0E",
    INIT_1c => x"ED204BCC1488ED5349CC1288ED444DCC1088ED4152CC016F846F46DE8E57F0BD",
    INIT_1d => x"01862188ED720ACC2688ED1F88ED0EC6BF861D88ED0101CC1B88ED0100CC1688",
    INIT_1e => x"8646DE8E57F0BD01C64F46DE8E5BF0BD03C64F2588A707862488A707862388A7",
    INIT_1f => x"206C616E7265746E6920676E69746F6F4208085BF07E01C64F01A7558684A7AA",
    INIT_20 => x"26FDD38C81EDA1EC34F48E10E5D38E6AF4BDEDF38E040A0D2E2E2E2E58454C46",
    INIT_21 => x"82F482F4C8DFC2DF82F476F400CD7EF7261EDE8C81EDA1EC4CF48E1000DE8EF7",
    INIT_22 => x"F07E9FF07E6CF07E63F07E5FF07E5BF07E57F07E72F46EF47AF482F47EF482F4",
    INIT_23 => x"9F6E08F89F6E04F89F6E06F89F6E0AF89F6E0CF89F6EC3F07EBFF07EA7F07EA3",
    INIT_24 => x"040A0D2E2E2E2064616F6C7075206B736944204D4F52206C61697265533900F8",
    INIT_25 => x"01C64F1EDEB700866AF4BD83F48E040A0D646564616F4C206B736944204D4F52",
    INIT_26 => x"E0260FC15C20DEF61FDEB626FC17F8265AC0A7EDF4BD5FFEFB1720DEF71FDEB7",
    INIT_27 => x"BD8435E0AB0434068D891F484848480E8D04346AF47EA0F48ED92630814C01C6",
    INIT_28 => x"B7038639018500E0B6390780EB2E1681EF2B11810A2F0981F72B3080FB2928F5",
    INIT_29 => x"DD8D0A2778850826018500E0B629DE7F28DE7F27DEB710863900E0B7118600E0",
    INIT_2a => x"00E0B6023439021A4FDC2627DE7AE12628DE7AE62629DE7A39021C01E0B6E620",
    INIT_2b => x"44204D4F52206D65646F6D580A0D3901E0B70235F120B38DF527788508260285",
    INIT_2c => x"550A0D046574656C706D6F432064616F6C70550A0D0464616F6C7055206B7369",
    INIT_2d => x"B7008625DEBF1AF68E23DEB70186B8FE1772F58E04726F7272452064616F6C70",
    INIT_2e => x"F61FDEB61FFB17F6265AC0A720252B00175FF9FA1720DEF71FDEB701C64F1EDE",
    INIT_2f => x"BE10346DFE169DF58E04FB176AF47E8BF58ED72630814C01C6DE260FC15C20DE",
    INIT_30 => x"F68E06260181903525DEBFED2684ADF1201AF68E4FFF1715860A2823FF1725DE",
    INIT_31 => x"8E062623DEB139FA1C39051A0326188139051A2EFF1706860826048139FA1C3A",
    INIT_32 => x"F68E24DEB7808621DE7FEF2623DEB14339FA1C1AF68E11FF17158639FA1C50F6",
    INIT_33 => x"072621DEB139041AFE1C7BF68E032624DE7A023521DEB721DEBB023439FA1C64",
    INIT_34 => x"4C080839FA1C1AF68EC4FE1715860435031F80C45A301F04340D20068623DE7C",
    INIT_35 => x"46042E4D4F5250206769666E6F63206D6F7266206B736964204D4F522064616F",
    INIT_36 => x"4D4F52040D0A2E2E2E6174616420676E6964616F6C202C434E595320646E756F",
    INIT_37 => x"756F4620746F4E206B736944204D4F52040D0A2E646564616F4C206B73694420",
    INIT_38 => x"00008C1F3015277C8D6C8D00008E20008E105A8D6AF4BD9DF68E040D0A2E646E",
    INIT_39 => x"F71FDEB701C61EDEB74F6AF4BDBFF68E6AF47EF0F68EEB2600008C101F31F326",
    INIT_3a => x"30814C01C6E1260FC15C20DEF61FDEB6ABF917F9265AC0A7678D5F82F91720DE",
    INIT_3b => x"BF46DFBFF92600008C1F3000008EC0E0B70086C0E0B702866AF47EDDF68EDA26",
    INIT_3c => x"FFCC46DF7947DF7948DF793949DF7844C0E0B6C0E0B70086C0E0B701863948DF",
    INIT_3d => x"B2FC17843549DFB6FB265ACE8D08C604343946DFB31055AACC072648DFB31000",
    INIT_3e => x"F4F78EF526F4F78C02300D2780E1E5F78E20C0022F60C1A5FC172086891F7F84",
    INIT_3f => x"000000040D0A3F2054414857ACF55806F750DDF246B2F44C0BF442946E87FC16"
    )

    port map (
	  do   => rdata0,
	  dop(0) => dp0,
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => wdata,
	  dip(0) => dp0,
	  en   => cs0,
	  ssr  => rst,
	  we   => we
	);

  ROM1 : RAMB16_S9
    generic map ( 
    INIT_00 => x"A780A610C6C0DF8E1074FE8E2EFA1AFB1EFB8FFBCEFCB9FC9BFCA1FC61F814F8",
    INIT_01 => x"17431FE4A7D0866AAFDD8C30FB265AE26F0CC65B0117E0DFBF00E08EF9265AA0",
    INIT_02 => x"0317A3FE8E0C0417F62A5A19048B0327856D0DC64FD0DF8E47031784FE8E9F04",
    INIT_03 => x"17408B981F5304175E86092C2081891FF1270D817F84370417B30217AAFE8E2E",
    INIT_04 => x"20F00217ACFE8EF52674FE8C02300F2780E13BFE8E20C0022F60C14704174C04",
    INIT_05 => x"17A4A60F0417A50317211F650217B2FE8E121F2D296B03173B341FBC2094ADC0",
    INIT_06 => x"27A4A1A4A7390F260D8117275E81DD271881E127088111285E0317070417A503",
    INIT_07 => x"0B031705201F30C0DF8E321FA20217BE203F31C2202131E503173F86E8031708",
    INIT_08 => x"279A03170527E4AC011FF0C4201F0634F0C41000C3101F390124E1AC20340629",
    INIT_09 => x"265A8E03172C031780A610C69603172E0317E4AEEE0117B2FE8E103439623203",
    INIT_0a => x"29B70217BC20EE265A7703172E8602237E810425208180A610C6E1AE860317F5",
    INIT_0b => x"3984A73F86A4AFA0A709273F8184A60F271035558DFFFF8E10341A24C0DF8C1E",
    INIT_0c => x"4AAF0427268D1F304AAE431F39FB265A188D08C6E3DF8E104603163F86490317",
    INIT_0d => x"A7A0A7A0A7FF8684A7A4A604263F8184A60A24C0DF8C21AEB9FE16480217068D",
    INIT_0e => x"0186398D46E0B7E086408D393D3139F7265A0427A1ACA0A608C6E3DF8E1039A0",
    INIT_0f => x"178D47E0B7208645E0B744E0B743E0B74F42E0B701862D8D47E0B7EF8641E0B7",
    INIT_10 => x"E0B6F926808547E0B63B341F4AAF00C08EF42600C28C80A740E0B6218D00C08E",
    INIT_11 => x"54545454A6E6D0DF8E104444444462A6363439F927088547E0B639F227408547",
    INIT_12 => x"FCBD8435FD265A20C60434B63562E762EA62A70F8462A65858585853A6E6E4E7",
    INIT_13 => x"0234A80117F12631813D273981230217F92653812A0217E2DF7F6802171186E3",
    INIT_14 => x"E0EB02340C2904358E01170434E46AE46AE4EBE0EBE0E6103421299101172629",
    INIT_15 => x"0117E26F1202161386E2DF731A02173F86BA27FFC102355FEB2080A70527E46A",
    INIT_16 => x"2320008310062762A3E4ECF901171286E3FCBDE4AF0130492562AC4D2930344A",
    INIT_17 => x"1780A684EB63EB62EB68011762AE750117981F03CB2F0017F3FE8E64E720C602",
    INIT_18 => x"10347120028D396532B701171486C326E4AC62AF5B0117981F53F526646A6501",
    INIT_19 => x"8D618D394AAF0229F68DF28D910017E50016F80016A101169035690017A4FE8E",
    INIT_1a => x"498D3944AF0229D58DD18D5E8D3946AF0229E08DDC8D728D3948AF0229EB8DE7",
    INIT_1b => x"8D3941A70229B18DB08D588D3942A70229BC8DBB8D6C8D3943A70229C78DC68D",
    INIT_1c => x"BF0016311FF48DB6FE8E39F726048180A63F011739C4A7808A0429A68DA58D5F",
    INIT_1d => x"8DC8FE8EE12044AED78DCEFE8EB4001643A6E18DD4FE8EF42048AEEA8DC2FE8E",
    INIT_1e => x"D02042A6B38DDFFE8ED92041A6BC8DDAFE8ECF204AAEC58DBCFE8ED82046AECE",
    INIT_1f => x"B2FE8EBF8DB88DB08DA98DA18D27FF17B2FE8E900016EBFE8EC4A6AA8DE4FE8E",
    INIT_20 => x"3C29088D011F42290E8DB800172D86121F4D29098DD520CE8DC78DC08D17FF17",
    INIT_21 => x"811D2530815B8D39E0AB04342829078D891F484848483229118D903561A71034",
    INIT_22 => x"3439021A39578003226681072561813937800322468112254181393080032239",
    INIT_23 => x"C602345120078B022F3981308B0F840235048D4444444402340235028D023510",
    INIT_24 => x"207F84048D0627E2DF7D00F09F6E8235F1265A3F8D438D2D860225E46880A608",
    INIT_25 => x"85E0DF9FA60234903501A6EE27018584A620E08E0926018584A6E0DFBE10342D",
    INIT_26 => x"3501A70235FA27028584A6E0DFBE1234458D2086008D8235018520E0B6052601",
    INIT_27 => x"A7FBDFFD0000CC30E08E39E2DFB7FF86016D84A7118684A70386E0DFBE138D90",
    INIT_28 => x"8D0427FEDF7D30E08E16345986028D1B86FEDF7F01E702C6FDDFFD04E703E702",
    INIT_29 => x"1A816C0027101B814100271008819635C5001784A70520098D042420810D2074",
    INIT_2a => x"51260A81110027100B812C0027100C81990027100D814500271016818E002710",
    INIT_2b => x"164A3327FBDFB67400165A3C0027105DFBDFFC9900168300261019C15CFBDFFC",
    INIT_2c => x"2710598116273DC1FEDFF65800160000CC5B00162500271050814CFBDFB66800",
    INIT_2d => x"2080FEDF7F39FDDFB70426FDDF7D39FEDF7F39FEDFB704263D81312754816E00",
    INIT_2e => x"A74C84E720C6FBDFB6168D0000CC1B20E12218C120C0FDDF7FFDDFF6ED224F81",
    INIT_2f => x"C15C4FF02650814CFBDFFC3903E702A7FBDFFDFCDFF64F39FEDF7FF726508102",
    INIT_30 => x"2650C15C84A702E7FBDFF72086FBDFF604E75F012519C15C04E6E78D5AEA2619",
    INIT_31 => x"FB0274FB0139FEDFF702E7FBDFF75FE4205F03E7FCDFF7082719C15CFCDFF6F4",
    INIT_32 => x"505EFA4CA5F847FDF8455CF94248FB1953FB183DFB1531FB105EFB047FFB0369",
    INIT_33 => x"94F9A7F8A7F8A7F8A7F894F992FC55D5F94488F958F1F853EDFB52A8F84DBCFA",
    INIT_34 => x"20204147504620524F4620342E312047554239305359530000000A0DFFFFFFFF",
    INIT_35 => x"43502020043D5053202004202D20043F54414857043E040000000A0D4B04202D",
    INIT_36 => x"20043D412020043D50442020043D58492020043D59492020043D53552020043D",
    INIT_37 => x"0000000000000000000004315343565A4E4948464504203A43432020043D4220",
    INIT_38 => x"300B2784AC1084AF1084EEAA558E10A0D08E84A7F086FB264A80A70F86F0FF8E",
    INIT_39 => x"2DA7D0DF8E10C0DFCE10FDFFB74444444443101F84EFD620ED26A0F08C00F089",
    INIT_3a => x"1084AF10AA558E1084EE2227A0F08C00F08930FB2A4AA66F0C862FA7F0862E6F",
    INIT_3b => x"2EA7D0DF8E10F186D520A5A70F88891F44444444101FD0DF8E1084EFE92684AC",
    INIT_3c => x"8EF32D0C814C80E7A66F0427A6E6211F4F2CE7A66F1420F92A4A0526A6E60C86",
    INIT_3d => x"9F6EC6DF9F6EC4DF9F6EC0DF9F6E62F816E2DFF753F9265A80A7A0A610C6F0FF",
    INIT_3e => x"0822CEDFBC8B300F27FFFF8CCCDFBE49584F4AAF80E64AAE431FCADF9F6EC8DF",
    INIT_3f => x"00FFB2FFC2FFBEFFBAFFB6FFC6FFB2FFC2DF9F6E42EE1F37F16E44AEC4EC1034"
    )

    port map (
	  do   => rdata1,
	  dop(0) => dp1,
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => wdata,
	  dip(0) => dp1,
	  en   => cs1,
	  ssr  => rst,
	  we   => we
	);

my_mon : process ( rw, addr, cs, rdata0, rdata1 )
begin
	 we    <= not rw;
	 case addr(11) is
	 when '0' =>
	   cs0   <= cs;
		cs1   <= '0';
		rdata <= rdata0;
    when '1' =>
	   cs0   <= '0';
		cs1   <= cs;
		rdata <= rdata1;
    when others =>
      null;
    end case;		
		
end process;

end architecture rtl;

