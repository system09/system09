    INIT_00 => x"D4C3FFC0BD45535255434552070346E46DE76EC2A7C4C2D3A7C4FFC0BD414552",
    INIT_01 => x"C600C843C98000AFC289C6E6C7D4C3FFC0BD4544494804060CE57EC0C8D413CD",
    INIT_02 => x"C01DC600C837C97FBCC289C6E6C7D4C3FFC0BD4C4145564552060629E87EC01D",
    INIT_03 => x"00C843C989C6F2C701BCC2B9C9D4C3FFC0BD4554414944454D4D490902D9E67E",
    INIT_04 => x"454C49504D4F435B09034BE67EC019E4C9E6FFC0BD5D275B0303C7E67EC01DC6",
    INIT_05 => x"C76FE37EE2D6C5FFC0BD454E4F5054534F50080362E57EC0C8D4C9E6FFC0BD5D",
    INIT_06 => x"4F54530506EEE67EC0C8D43500DCC2B3C5D5E3E6D4E6D4D5E87BC29EC8BAE6E6",
    INIT_07 => x"1BBCC20CC2DBC7FDE87BC2D4C8F2C7D6C50CC2DBC7AFC0E6C7F7C1FFC0BD3F50",
    INIT_08 => x"E804D5FCC066E7FFC0BD3A0102ADE87EC0E2C8D6C530E637C9E4BCC2D4C8F2C7",
    INIT_09 => x"DB42CCFCC0AFC2A7C4FFC0BD454D414E4F4E3A070217E77EC0BFCDCCC5BFC52E",
    INIT_0a => x"E6C766E7FFC0BD544E4154534E4F43080201E77EC0D5E3BFCDCCC5CCC504D56A",
    INIT_0b => x"52415608022CE97EC0FDCC3AC17EC0E8CC4FC173E97BC289CD80BCC28000AFC2",
    INIT_0c => x"66E7FFC0BD45554C4156050211E47EC0DACCB3C525C166E7FFC0BD454C424149",
    INIT_0d => x"97E87EC0B4C6AEC9D5C0BDEEC0BD474E495254534F44080414E97EC0E8CC63C1",
    INIT_0e => x"CCC5FDCCE6C76DC801BCC237C9FF00AFC2B2E966E7FFC0BD474E495254530606",
    INIT_0f => x"DDC67EC889C6D1C6AEC9E6C727C2FFC0BD2928244F54050446E87EC0DACCFDCC",
    INIT_10 => x"C989C60BC789C6D1C6AEC9E6C727C2FFC0BD2928244F542B0604FEE77EC0C2D3",
    INIT_11 => x"29282452434E49070464E87EC0A2D363C6DDC6E6C700C8D7C9B4C60BC77EC8E0",
    INIT_12 => x"C21DC6D7C9B4C60BC768EA7BC21BC989C60BC789C6D1C6AEC9E6C727C2FFC0BD",
    INIT_13 => x"DCC2CBC263C170EA40EA0EEAEFE9B2E900007EC02BC7DBC77EC063C6DDC601BC",
    INIT_14 => x"03047CE97EC02700CBC2A7C4E8CCC5C3FFC0BD5453494C584650070413E8F0C2",
    INIT_15 => x"42C8D0EA7BC2D4C895C654C7C5C36CCC95C650CCE6C742CCC9E6FFC0BD584650",
    INIT_16 => x"E907D3E0BCC2B4EA98C2E6C795C650CC7EC0E8CCE8CC42D595C6D7C91FC826CC",
    INIT_17 => x"7EC0A3EA02BCC2FFC0BD4F542B0307DCE87EC0A3EA00BCC2FFC0BD4F540203E9",
    INIT_18 => x"BD53454C424149524156090685EA7EC0A3EA04BCC2FFC0BD52434E49040787E8",
    INIT_19 => x"A7C4C3C6DDC6ACD4FFC0BD455355463C0504E2EA7EC0A2C1DACC7ACC66E7FFC0",
    INIT_1a => x"C2E8CCC3C626CCDACCFEBCC263EB7BC237C90EC9B9C9A7C428C4D4C895C650CC",
    INIT_1b => x"C092C0ABC835EBFFC0BD544958453F0507D3E57EC0D1C626CCE8CCC3C669EB6E",
    INIT_1c => x"C0BFCD01BCC2E8CCE6C7A7C498C27BC2ABC835EBFFC0BD4649020303EB7EC0AF",
    INIT_1d => x"C0BD454C4948570503F2EA94EB6EC26EC2E6D4FFC0BD4441454841050386EB7E",
    INIT_1e => x"A7C495D401BCC2D3CDACD4FFC0BD4E454854040395E97EC012CE01BCC289EBFF",
    INIT_1f => x"C0D5E3BFCD02BCC2A7C4ACD4FFC0BD4E494745420503A9E97EC0D5E32CC600C8",
    INIT_20 => x"7EC0E8CC98C27BC2ABC835EB95D402BCC2D3CDFFC0BD4C49544E550503B8EB7E",
    INIT_21 => x"450403B3E67EC0E8CC6EC2E6D495D402BCC2D3CDFFC0BD4E49414741050304EC",
    INIT_22 => x"29ECFFC0BD54414550455206032FEB7EC0D2EB12CE01BCC2AAEBFFC0BD45534C",
    INIT_23 => x"A4EB7EC0BFCD03BCC2E8CCE6C7A7C407C3E6D4FFC0BD4F44020354EC7EC0D2EB",
    INIT_24 => x"03BCC2D3CDFFC0BD504F4F4C04039FEA71EC6EC225C3E6D4FFC0BD4F443F0303",
    INIT_25 => x"FFC0BD504F4F4C2B05033EEC7EC02CC600C8A7C4E8CC26CCE6C73DC3E6D495D4",
    INIT_26 => x"EC7BC295D4CCC5D3CDFFC0BD3B010323ECA6EC6EC262C3E6D495D403BCC2D3CD",
    INIT_27 => x"5202074FE77EC0D2EB7EC0E6D4FFC0BD7D010770EB7EC0F4D47EC0E6D44DE8E3",
    INIT_28 => x"ABC835EBFFC0BD45523F0307D2EC7EC0E8CC42CC13CDD4C36EC2E6D4FFC0BD45",
    INIT_29 => x"4E4F4F4406042AE67EC0D2EB01EDFFC0BD7D4552030715EB08ED6EC27BC298C2",
    INIT_2a => x"A1E47EC01DC62D00CBC2E6C7B9C91DC654C7B9C95BC589C6D5C0BDEEC0BD594C",
    INIT_2b => x"45EDBD594C4E4F040281EC7EC01DC6F0C389C6D5C0BDEEC0BD434F564F440504",
    INIT_2c => x"046AEDBD454449534E49060050E980ED026AEDBD4854524F46050067EC000000",
    INIT_2d => x"EDBD52454C424D45535341090007EA9FED066AEDBD41525458450500EEEC8FED",
    INIT_2e => x"D7C902BCC289C6E6C7A7C3A7C4FFC0BD5453494C44524F570802B7ECAEED086A",
    INIT_2f => x"C80EC9F0C34CC5FFC0BD4F534C410400C7ED7EC089C62300CBC2E6C7E8CCFDCC",
    INIT_30 => x"455250080061ED7EC01DC6F0C32D00DCC2FFBCC289C6F0C330E637C9CFBCC2AB",
    INIT_31 => x"ED7EC02D00F0C230E637C9CEBCC2ABC80EC95BC5AEC9F0C3FFC0BD53554F4956",
    INIT_32 => x"470B00A5ED7EC01DC65BC589C6F0C3FFC0BD534E4F4954494E494645440B003B",
    INIT_33 => x"45525255432D5445530B0038EA7EC089C65BC5FFC0BD544E45525255432D5445",
    INIT_34 => x"C889C654C7A7C3FFC0BD454D414E434F560704FEEC7EC01DC65BC5FFC0BD544E",
    INIT_35 => x"46C79BEE98C2E6C795C6AEC97EC037C91FBCC2B4C628CD6CCC42C8B4EE7BC2D4",
    INIT_36 => x"524544524F0500F1ED7EC0B0CF96EEFFC0BD434F562E0406CDEB7EC03F017DD5",
    INIT_37 => x"8DD5F4EE3DC37BCFCEEEB4C6FEEE07C300BCC2E0C9F2C75BC5F0C3ECE0FFC0BD",
    INIT_38 => x"C0F6ED8CEDF6EDABED7DEDFFC0BD4853455246050086ED7EC0CEEE89C6203A02",
    INIT_39 => x"0704DAEE7EC067EDDBC7D0ED66E7FFC0BD5952414C554241434F560A0693EC7E",
    INIT_3a => x"8FC8E0C93AC595C688C366EF07C303BCC223BCC2CCC5FFC0BD41464E504F5421",
    INIT_3b => x"D1C6FFC0BD4C494154525543070476EE7EC02900CBC2D7C93AC556EF62C3B3C5",
    INIT_3c => x"524F4628070424EF7EC02BC784EF98C289CD75C7E6C795C6D7C90BC78AEF6EC2",
    INIT_3d => x"C52CC688C37BEFFDBCC295C688C3C5EF07C303BCC223BCC2A7C4FFC0BD544547",
    INIT_3e => x"FEBCC2C5C32500CBC27BEF02BCC2B6C32300CBC27BEF01BCC2A7C3B2EF62C3B3",
    INIT_3f => x"C67EE2D6C5FFC0BD544547524F4606021CEE7EC047EFDACCE0C92700CBC27BEF",
