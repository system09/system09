    INIT_00 => x"0EC9F2C7A7C4E0C937C902BCC265CD00C896CCE6C728CDBAE699E389C65BC5B4",
    INIT_01 => x"8000AFC289C6D4C3FFC0BD45564F4D455206068EEE7EC0A3EF30E637C9F1BCC2",
    INIT_02 => x"52454B52414D4F4408042EF00BF06EC27BCFB0CFB4C6E6C7D4C34DE8AFC037C9",
    INIT_03 => x"A2D3AEC9E0C9F2C75BC52D00CBC2E6C7B4C626CCA3EF95C6E6C7D5C0BDEEC0BD",
    INIT_04 => x"C5A7C4FDCCE6C7F0C3E8CC60F066E7A7C4FFC0BD52454B52414D0602B4ED7EC0",
    INIT_05 => x"D1C695C6BFC4FFC0BD57454E4104063FEF7EC0A2D3DACCE6C7AEC9E0C9F0C35B",
    INIT_06 => x"C9E6C7F5F07BC2C9C737C9F2C86FE330E637C9E0BCC2ABC889C6E6C7D9D3D6C5",
    INIT_07 => x"EE7EC08CF02CC6BFC4DDC670C0F5F07BC2C9C737C9D4C860F0AFC26CCC95C6AE",
    INIT_08 => x"95C682C44300DCC20008AFC24300CBC200F8AFC2FFC0BD4D454D49482106045E",
    INIT_09 => x"0602C1E97EC014F17BC2E2C860C92CC682C4F2C795C682C42CC682C460C9E6C7",
    INIT_0a => x"1F4F444C4F43040695ED7EC0E0C9A7C4E0C920BCC282C4FFC0BD444553554E55",
    INIT_0b => x"CBC200BCC247EF09F19ACB65BCC200BCC23AC5FFC0BDFE01CE06357E01CE108B",
    INIT_0c => x"7279706F431F8DD559CF54E100BCC259CFE4C17FBCC24EEE12EFDBC71DD52F00",
    INIT_0d => x"531D8DD559CF67672D6874726F46204343482035303032202963282074686769",
    INIT_0e => x"82C459CF72656E6265754820736E61482079622074726F702039306D65747379",
    INIT_0f => x"442806049BEFFAE559CF59CF4D415220426B20078DD53CD209BCC288C90ABCC2",
    INIT_10 => x"D4F2C7CCC5D3CDFFC0BD3E53454F440503FDF17EC03DCDDDC6FFC0BD3E53454F",
    INIT_11 => x"BCC266E7FFC0BD45444F43040215ED7EC0D5E36ADBD5C0AFC204F2E6D4BFCD95",
    INIT_12 => x"CCC5D3CDFFC0BD45444F433B05033FF17EC0BFCD05BCC2BFC52EE8BEEDDACCFD",
    INIT_13 => x"C016E9FFC0BD3A52454F4405062BED7EC0F4D4BEED04F2E6D4BFCD05BCC295D4",
    INIT_14 => x"C0DACC03BCC239F2FFC0BD45444F4352454F44080642EE7EC06ADBD5C0AFC2EB",
    INIT_15 => x"EE4DE8BFF27BC295D405BCC2D3CDFFC0BD45444F432D444E450808B2F07EC0EB",
    INIT_16 => x"414E45060673EF7EC02CC6AEC9FFC0BD524F5443455621070634F27EC0F6ED25",
    INIT_17 => x"3BBCC2FFC0BD454C424153494407060CEF7EC01DC600C87EBCC2FFC0BD454C42",
    INIT_18 => x"EF7EC02CC6BFC437C9E2E895C6BFC4FFC0BD594E414D0406A6F27EC01DC600C8",
    INIT_19 => x"43C9E2E8D4C80BC73700CBC200BCC2D1C6AEC937C4FFC0BD53454D49540506F1",
    INIT_1a => x"5344524F570B0409F37EC02CC6BFC400BCC23700CBC2DDC67EC02BC748F37BC2",
    INIT_1b => x"C2D4C876CD54C783F37BC2E6C795C696CC71F36EC200C8FFC0BD52455050494B",
    INIT_1c => x"C7D7C924BCC25CC43CC61DD5FFC0BD5344524F5728060422F37EC042C86FF37B",
    INIT_1d => x"88C370C0A1C65CC488C3C8F307C354C79ACB20BCC2F2C703BCC2E0C920BCC2E6",
    INIT_1e => x"7BC295C688C304F407C375C7FFBCC2CCC5D1C600BCC259CFB6F362C3B3C52CC6",
    INIT_1f => x"B3C588C3E0C93AC595C688C346C7FEF37BC20EC9E0C93AC595C688C3F2C7FEF3",
    INIT_20 => x"C03CD200BCC2ECE0DDC659CF46C7DBC721F47BC243C9E2E846CE42C8DAF362C3",
    INIT_21 => x"BCC2E6C7B4C6E6C795C6E6C7D1C6AEC9DDC659CF2EF47BC20EC968C43CBCC27E",
    INIT_22 => x"C65CC496CC7BCFB0CF48CF7EBCC237C91FBCC255F46EC2D6C54DF47BC228C920",
    INIT_23 => x"F366F3AFC289C6F0C3FFC0BD5344524F57050053F2CFF36EC22CC600C870C0A1",
    INIT_24 => x"EBEB7EC091F370C0AFC295C6AFC2FFC0BD5344524F574C4C410806DCF27EC091",
    INIT_25 => x"44412E0404A1F47EC01DC65CC442C873D146CEFF00AFC2FFC0BD21522E580404",
    INIT_26 => x"3CD289C65CC4FFC0BD455459422E050457F07EC026D2C4C989C65CC4FFC0BD52",
    INIT_27 => x"74F27EC048CF6DC8D6C537C928C97FBCC2E6C7FFC0BD4353412E0404C9EE7EC0",
    INIT_28 => x"C921F57BC228C906BCC2E6C75DC810BCC295C6CCC4A6F4FFC0BD504D55440402",
    INIT_29 => x"D7C988C3E6C74AF507C300BCC20BC77BCFC1F459CFE6C700C8D7C9F2C7D1C6C4",
    INIT_2a => x"D557F53DC3EAF4B4C65FF507C300BCC20BC77C018DD53AF53DC37BCFD7F489C6",
    INIT_2b => x"0504C8F27EC02BC746C729F57BC243C9E2E80EC90BC7E0C900C854C7207C028D",
    INIT_2c => x"E6C7B9C900C837C989CDA7C43AC5F2C70EC9F2C70003AFC2FFC0BD3F3F414643",
    INIT_2d => x"C789C6F2C7DDC6B9C9D1C601BCC2AFC0E6C737C937C989CD7FBCC221BCC289C6",
    INIT_2e => x"C9F2C7D6C5AEC9E5F57BC289CD7FBCC221BCC27EC0F2C846C7CDF57BC2D4C854",
    INIT_2f => x"AFC0E6C737C985F5E6C7FFC0BD3F414643040478ED7EC0CCC546C7B5F57BC237",
    INIT_30 => x"B9C922F698C2E6C795C696CCAFC0E6C737C9ABC828C976CDF2C789C6A7C328CD",
    INIT_31 => x"F2F27EC0CCC5DBC77EC085F513CD38F67BC289CD20BCC200BCC289C6E6C77EC0",
    INIT_32 => x"CFB4C628CDB0CF18C7EAC620202D2D2020067DD5E6C7FFC0BD444145482E0504",
    INIT_33 => x"CD2072656F64058DD5E6C785F67BC2F3F5E6C76CCC95C6AEC9E6C7B0CF18C7B0",
    INIT_34 => x"2E0604BCF47EC064726F5720058DD5CEEE76CD28CDB0CFFBC6DBC7B0CFB4C628",
    INIT_35 => x"B0CFB4C628CD8ECFD7C904BCC2C4C9C4C937C901BCC2F2C7FFC0BD4E454B4F54",
    INIT_36 => x"F4E6C7B4C6E6C7203A028DD5C1F4E6C759CFFFC0BD4D4F43454405049EF67EC0",
    INIT_37 => x"01BCC2F2C7D6C5C1F495C6E6C77BCFEAF47BCFD7F4E6C789C67BCFEAF47BCFD7",
    INIT_38 => x"C77EC0AEC947F6E6C71FF77BC2F3F5E6C77BCF48CFD7C90EBCC20BF77BC237C9",
    INIT_39 => x"C992C0F3F595C6E6C792C0F3F5E6C7AEC9A5F695C6E6C743F77BC2F3F595C6E6",
    INIT_3a => x"7EC0DBC754F77BC2E2E8CBF6A6F4FFC0BD4545534D040686F47EC0AEC97EC0AE",
    INIT_3b => x"BDEEC0BD4553414246464F4408048CF27EC04FF7C9E6FFC0BD45455303026EF4",
    INIT_3c => x"30E62CC6CCC4DDC6F2D290E5AFC27EE2D6C52CC6CCC489C6D1C695C6CCC4D5C0",
    INIT_3d => x"BD58480201D1F47EC06EE8FDCC7CF766E7FFC0BD455341424646060401F57EC0",
    INIT_3e => x"4E4548545B06017FF5027FF7BD4E420201C6F70A7FF7BD4D4402018AF3107FF7",
    INIT_3f => x"DBC700F86EC2FFC0BD5D4C414E4F495449444E4F435B0D0463F77EC0FFC0BD5D",
