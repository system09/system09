--
-- Ram1k_b4.vhd
--
-- 1K Byte RAM made out of 2 x 512 byte Block RAMs.
-- John Kent
-- 3 February 2007
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
library unisim;
	use unisim.vcomponents.all;

entity ram1k is
    Port (
       WB_CLK_I : in  std_logic;
       WB_RST_I : in  std_logic;
       WB_ADR_I : in  std_logic_vector (9 downto 0);
       WB_DAT_O : out std_logic_vector (7 downto 0)
       WB_DAT_I : in  std_logic_vector (7 downto 0);
       WB_WE_I  : in  std_logic;
       WB_STB_I : in  std_logic;
    );
end ram1k;

architecture rtl of ram_2k is

   signal rdata0   : std_logic_vector (7 downto 0);
   signal rdata1   : std_logic_vector (7 downto 0);
   signal ena0     : std_logic;
   signal ena1     : std_logic;

   component RAMB4_S8
    generic (
      INIT_00, INIT_01, INIT_02, INIT_03,
      INIT_04, INIT_05, INIT_06, INIT_07,
      INIT_08, INIT_09, INIT_0A, INIT_0B,
      INIT_0C, INIT_0D, INIT_0E, INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
    );

    port (
      clk, we, en, rst : in std_logic;
      addr :  in std_logic_vector(8 downto 0);
      di   :  in std_logic_vector(7 downto 0);
      do   : out std_logic_vector(7 downto 0)
    );
  end component;

begin

  MY_RAM0 : RAMB4_S8
    generic map ( 
INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000", INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000"    )

    port map ( 
	clk => WB_CLK_I,
	en  => ena0,
	we  => WB_WE_I,
	rst => WB_RST_I,
	addr(8 downto 0) => WB_ADR_I(8 downto 0),
	di(7 downto 0)   => WB_DAT_I(7 downto 0),
	do(7 downto 0)   => rdata0(7 downto 0)
	);

  MY_RAM1 : RAMB4_S8
    generic map ( 
INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000", INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000"    )

    port map ( clk => clk,
	clk => WB_CLK_I,
	en  => ena1,
	we  => WB_WE_I,
	rst => WB_RST_I,
	addr(8 downto 0) => WB_ADR_I(8 downto 0),
	di(7 downto 0)   => WB_DAT_I(7 downto 0),
	do(7 downto 0)   => rdata1(7 downto 0)
	);


my_ram_1k : process (WB_STB_I, WB_ADR_I, rdata0, rdata1 )
begin
	case WB_ADR_I(9) is
	when "0" =>
		ena0     <= WB_STB_I;
		ena1     <= '0';
		WB_DAT_O <= rdata0;
	when "1" =>
		ena0     <= '0';
		ena1     <= WB_STB_I;
		WB_DAT_O <= rdata1;
	when others =>
		null;
	end case;

end process;

end;

