--===========================================================================--
--                                                                           --
--  dpr_2k.vhd - Synthesizable 2KB Dual Port RAM using Xilinx 18KBit BLKRAM  --
--                                                                           --
--===========================================================================--
--
--  File name      : dpr_2k.vhd
--
--  Purpose        : Implement 2KByte Dual Port RAM
--
--  Dependencies   : ieee.std_logic_1164
--                   ieee.std_logic_arith
--                   unisim.vcomponents
--
--  Author         : John E. Kent
--
--  Email          : dilbert57@opencores.org      
--
--  Web            : http://opencores.org/project,system09
--
--  dpr_2k.vhd 2KByte Dual Port Block RAM Instantiation written in VHDL.
-- 
--  Copyright (C) 2010 John Kent
--
--  This program is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
--===========================================================================--
--                                                                           --
--                              Revision  History                            --
--                                                                           --
--===========================================================================--
--
-- Version Author        Date           Changes
-- 0.1     John Kent     7th June 2010  Added header & GPL
--
library IEEE;
   use ieee.std_logic_1164.all;
   use ieee.std_logic_arith.all;

library unisim;
	use unisim.vcomponents.all;

entity dpr_2k is
    Port (
       --
       -- Port A
       --
       clk_a      : in  std_logic;
       rst_a      : in  std_logic;
       cs_a       : in  std_logic;
       rw_a       : in  std_logic;
       addr_a     : in  std_logic_vector (10 downto 0);
       data_in_a  : in  std_logic_vector (7 downto 0);
       data_out_a : out std_logic_vector (7 downto 0);
       --
       -- Port B
       --
       clk_b      : in  std_logic;
       rst_b      : in  std_logic;
       cs_b       : in  std_logic;
       rw_b       : in  std_logic;
       addr_b     : in  std_logic_vector (10 downto 0);
       data_in_b  : in  std_logic_vector (7 downto 0);
       data_out_b : out std_logic_vector (7 downto 0)
    );
end entity;

architecture rtl of dpr_2k is


signal we_a : std_logic;
signal dp_a : std_logic_vector(0 downto 0);
signal we_b : std_logic;
signal dp_b : std_logic_vector(0 downto 0);

begin

  ROM : RAMB16_S9_S9
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map (
	  doa     => data_out_a,
	  dopa    => dp_a,
	  addra   => addr_a,
	  clka    => clk_a,
	  dia     => data_in_a,
	  dipa    => dp_a,
	  ena     => cs_a,
	  ssra    => rst_a,
	  wea     => we_a,
	  dob     => data_out_b,
	  dopb    => dp_b,
	  addrb   => addr_b,
	  clkb    => clk_b,
	  dib     => data_in_b,
	  dipb    => dp_b,
	  enb     => cs_b,
	  ssrb    => rst_b,
	  web     => we_b
	);

my_ram_2k : process ( rw_a, rw_b )
begin
  we_a    <= not rw_a;
  we_b    <= not rw_b;
end process;

end architecture;

