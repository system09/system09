library IEEE;
   use IEEE.std_logic_1164.all;
   use IEEE.std_logic_arith.all;
library unisim;
   use unisim.vcomponents.all;

entity SYS09BUG_F000 is
   port(
      clk    : in  std_logic;
      rst    : in  std_logic;
      cs     : in  std_logic;
      rw     : in  std_logic;
      addr   : in  std_logic_vector(10 downto 0);
      rdata  : out std_logic_vector(7 downto 0);
      wdata  : in  std_logic_vector(7 downto 0)
   );
end SYS09BUG_F000;

architecture rtl of SYS09BUG_F000 is

   type data_array is array(0 to 3) of std_logic_vector(7 downto 0);
   signal xdata : data_array;
   signal en : std_logic_vector(3 downto 0);
   signal we : std_logic;

component RAMB4_S8
generic (
   INIT_00, INIT_01, INIT_02, INIT_03,
   INIT_04, INIT_05, INIT_06, INIT_07,
   INIT_08, INIT_09, INIT_0A, INIT_0B,
   INIT_0C, INIT_0D, INIT_0E, INIT_0F : bit_vector (255 downto 0)
    );
   port (
      clk, we, en, rst : in std_logic;
      addr : in std_logic_vector(8 downto 0);
      di   : in std_logic_vector(7 downto 0);
      do   : out std_logic_vector(7 downto 0)
      );
     end component RAMB4_S8;

   begin

   ROM00: RAMB4_S8
      generic map (
         INIT_00 => x"8C02300D2780E12CF08E20C0022F60C10AF89FAD2086891F7F8406F89FAD02F0",
         INIT_01 => x"CD8E040D0A3F2054414857BCF258EAF0463EF042946E29021635F08EF52635F0",
         INIT_02 => x"B6B035EE261F30F6263F310A254700E0B6E2048E10E8038E30343B341F4AAF00",
         INIT_03 => x"0235ED261F30F5263F310C25474700E0B6E2048E10E8038E02343034B03501E0",
         INIT_04 => x"2E2E2E6B7369642045444920676E6974616D726F460D0AB03501E0B70235B035",
         INIT_05 => x"6E20657669726420454449040D0A043F207265626D754E2065766972440D0A20",
         INIT_06 => x"6574656C706D6F432074616D726F460D0A04202164657461636F6C6C6120746F",
         INIT_07 => x"002510308169FF17FB2450FF1753F2BD89F08EBDF4BD04204B53494445444904",
         INIT_08 => x"017FFB265A80A75F4F00028E3AF5BDFD008E0001F7891F3080E90022103381EF",
         INIT_09 => x"F60101B601A70186846C042600814C0201B684A70101B600028E0201B7018601",
         INIT_0a => x"028EC82600810101B601017C0201B70186D72600810201B602017C15F5BD0201",
         INIT_0b => x"8EF1F4BDFFC64F00028E15F5BDFFC6FF86016F846F00028EF1F4BDFFC6FF8600",
         INIT_0c => x"8E102034016F846F00028EF1F4BD03C64F00028E15F5BDFFC64F016F846F0002",
         INIT_0d => x"FFC6FF861D88ED0101CC1B88ED0001F64F2035F72618C15C85A7A0A610C6E1F0",
         INIT_0e => x"F5BD03C64F2588A707862488A707862388A701862188ED01FECC2688ED1F88ED",
         INIT_0f => x"E0B7038639018500E0B653F27ECFF08E2503170201F70101B701C64F00F78E15"
      )
      port map (
         clk     => clk,
         en      => en(0),
         we      => we,
         rst     => rst,
         addr    => addr(8 downto 0),
         di      => wdata,
         do      => xdata(0)
      );

   ROM01: RAMB4_S8
      generic map (
         INIT_00 => x"20DD8D0A2778850826018500E0B60A017F09017F0801B710863900E0B7118600",
         INIT_01 => x"8500E0B6023439021A4FDC2608017AE12609017AE6260A017A39FD1C01E0B6E6",
         INIT_02 => x"646F6D580A0D39F826048180A6E78D3901E0B70235F120B38DF5277885082602",
         INIT_03 => x"706D6F432064616F6C70550A0D0464616F6C7055206B73694420454449206D65",
         INIT_04 => x"626D754E2065766972440A0D04726F7272452064616F6C70550A0D046574656C",
         INIT_05 => x"175AF28E04294E2F5928203F206572755320756F59206572410A0D043A207265",
         INIT_06 => x"01B730802801221033812E01251030816AFF17FB293CFF178BFF1794F28E91FF",
         INIT_07 => x"815F843DFF17FB290FFF175EFF17A5F28E4BFF17308B0001B66CFF1794F28E00",
         INIT_08 => x"0101B701C64F00028E0401B701860601FF2DF4CEB10117B3265981FF0027104E",
         INIT_09 => x"D501170201F60101B600028ED6002510E00017870117E0002510EA00170201F7",
         INIT_0a => x"B00017570117B0002510BA00170201F70101B75C0201F60101B600028E710117",
         INIT_0b => x"0101B75C0201F60101B600028E410117A501170201F60101B600028EA6002510",
         INIT_0c => x"88E60B01B74C2688A600028E76002510800017270117800025108A00170201F7",
         INIT_0d => x"01F70101B700028E5C0201F60101B60301176701170201F60101B60C01F75C27",
         INIT_0e => x"00173701170201F60101B600028E38002510420017E90017420025104C001702",
         INIT_0f => x"01F70101B701C64F00F78EC3260B01B14C01C6CB260C01F15C0201F60101B6D3"
      )
      port map (
         clk     => clk,
         en      => en(1),
         we      => we,
         rst     => rst,
         addr    => addr(8 downto 0),
         di      => wdata,
         do      => xdata(1)
      );

   ROM02: RAMB4_S8
      generic map (
         INIT_00 => x"CE1BFE1715860A28EFFD170601FE403443FE1685F28E53F27E73F28E11011702",
         INIT_01 => x"FAFD1706860826048139FA1C4DF4CE06260181C0350601FFED26C4ADF1202DF4",
         INIT_02 => x"2DF4CEDDFD17158639FA1C63F4CE06260401B139FA1C39051A0326188139051A",
         INIT_03 => x"350301B70301BB023439FA1C77F4CE0501B7808603017FEF260401B14339FA1C",
         INIT_04 => x"043439041AFE1C2DF4CE04017C0B260301B139FA1C80A78EF4CE032605017A02",
         INIT_05 => x"0600CC82357FFD170686023439FA1C2DF4CE8CFD1715860435011F80C45A101F",
         INIT_06 => x"E4E606E1FD5A4F023401C64F668DD602160CE1FDE000CC1EE1FD0200CC1EE1FD",
         INIT_07 => x"8E102034AC02170EE1FD2000CCE48D82355F04E1FD01C60AE1FD0001F608E1FD",
         INIT_08 => x"8802170EE1FD3000CCC08D395F9502172035F4263F3180E700E1FCB202170001",
         INIT_09 => x"0123038103A6395F7002172035F4263F3100E1FD80E68D02174F00018E102034",
         INIT_0a => x"00000000000000000000000000000000000000000000395F03A6395F0001B74F",
         INIT_0b => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0c => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0d => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0e => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0f => x"0000000000000000000000000000000000000000000000000000000000000000"
      )
      port map (
         clk     => clk,
         en      => en(2),
         we      => we,
         rst     => rst,
         addr    => addr(8 downto 0),
         di      => wdata,
         do      => xdata(2)
      );

   ROM03: RAMB4_S8
      generic map (
         INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_08 => x"270281358D00C48E1000C3FDF18CECFFC0CE1000000000C00000000000000B20",
         INIT_09 => x"5D891F158DD08CA71A8DD48CA71F8DEA20DA8CA7268DDE8CA72B8DF626168110",
         INIT_0a => x"8D0B2784EC00C38E0F2600C48C10C920F5265A80A71435098D1434C58CAED927",
         INIT_0b => x"C60AE1FD908CE608E1FDE4E606E1FD5A4F02349B9C6E39A0A604C38E109D2626",
         INIT_0c => x"3F3180E700E1FC1E8D00018E102034178D0EE1FD2000CCE48D82355F04E1FD01",
         INIT_0d => x"0039F92708C50EE1FC39F22740C50EE1FCF92680C50EE1FC395F028D2035F526",
         INIT_0e => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_0f => x"0000000000000000000000000000000000000000000000000000000000000000"
      )
      port map (
         clk     => clk,
         en      => en(3),
         we      => we,
         rst     => rst,
         addr    => addr(8 downto 0),
         di      => wdata,
         do      => xdata(3)
      );

   rom_glue: process (cs, rw, addr, xdata)
   begin
      en <= (others=>'0');
      case addr(10 downto 9) is
      when "00" =>
         en(0)  <= cs;
         rdata  <= xdata(0);
      when "01" =>
         en(1)  <= cs;
         rdata  <= xdata(1);
      when "10" =>
         en(2)  <= cs;
         rdata  <= xdata(2);
      when "11" =>
         en(3)  <= cs;
         rdata  <= xdata(3);
      when others =>
         null;
      end case;
      we <= not rw;
   end process;
end architecture rtl;

library IEEE;
   use IEEE.std_logic_1164.all;
   use IEEE.std_logic_arith.all;
library unisim;
   use unisim.vcomponents.all;

entity SYS09BUG_F800 is
   port(
      clk    : in  std_logic;
      rst    : in  std_logic;
      cs     : in  std_logic;
      rw     : in  std_logic;
      addr   : in  std_logic_vector(10 downto 0);
      rdata  : out std_logic_vector(7 downto 0);
      wdata  : in  std_logic_vector(7 downto 0)
   );
end SYS09BUG_F800;

architecture rtl of SYS09BUG_F800 is

   type data_array is array(0 to 3) of std_logic_vector(7 downto 0);
   signal xdata : data_array;
   signal en : std_logic_vector(3 downto 0);
   signal we : std_logic;

component RAMB4_S8
generic (
   INIT_00, INIT_01, INIT_02, INIT_03,
   INIT_04, INIT_05, INIT_06, INIT_07,
   INIT_08, INIT_09, INIT_0A, INIT_0B,
   INIT_0C, INIT_0D, INIT_0E, INIT_0F : bit_vector (255 downto 0)
    );
   port (
      clk, we, en, rst : in std_logic;
      addr : in std_logic_vector(8 downto 0);
      di   : in std_logic_vector(7 downto 0);
      do   : out std_logic_vector(7 downto 0)
      );
     end component RAMB4_S8;

   begin

   ROM00: RAMB4_S8
      generic map (
         INIT_00 => x"A780A610C6C0DF8E1074FE8E2EFA1AFB1EFB8FFBE0FCC5FC9BFCA1FC61F814F8",
         INIT_01 => x"17431FE4A7D0866AAFDD8C30FB265AE26F0CC65B0117E0DFBF00E08EF9265AA0",
         INIT_02 => x"0317A3FE8E0C0417F62A5A19048B0327856D0DC64FD0DF8E47031784FE8EB504",
         INIT_03 => x"17408B981F6504175E86092C2081891FF1270D817F84370417B30217AAFE8E2E",
         INIT_04 => x"20F00217ACFE8EF52674FE8C02300F2780E13BFE8E20C0022F60C15904175E04",
         INIT_05 => x"17A4A6210417A50317211F650217B2FE8E121F2D296B03173B341FBC2094ADC0",
         INIT_06 => x"27A4A1A4A7390F260D8117275E81DD271881E127088111285E0317190417A503",
         INIT_07 => x"0B031705201F30C0DF8E321FA20217BE203F31C2202131F703173F86FA031708",
         INIT_08 => x"27A603170527E4AC011FF0C4201F0634F0C41000C3101F390124E1AC20340629",
         INIT_09 => x"265AA003172C031780A610C6A803172E0317E4AEEE0117B2FE8E103439623203",
         INIT_0a => x"29B70217BC20EE265A8903172E8602237E810425208180A610C6E1AE980317F5",
         INIT_0b => x"3984A73F86A4AFA0A709273F8184A60F271035558DFFFF8E10341A24C0DF8C1E",
         INIT_0c => x"4AAF0427268D1F304AAE431F39FB265A188D08C6E3DF8E105803163F865B0317",
         INIT_0d => x"A7A0A7A0A7FF8684A7A4A604263F8184A60A24C0DF8C21AEB9FE16480217068D",
         INIT_0e => x"E1FD0200CC1EE1FD0600CC393D3139F7265A0427A1ACA0A608C6E3DF8E1039A0",
         INIT_0f => x"178D0EE1FD20C60AE1FD08E1FD06E1FD5F04E1FD0100CC2E8D0CE1FDE000CC1E"
      )
      port map (
         clk     => clk,
         en      => en(0),
         we      => we,
         rst     => rst,
         addr    => addr(8 downto 0),
         di      => wdata,
         do      => xdata(0)
      );

   ROM01: RAMB4_S8
      generic map (
         INIT_00 => x"E1FCF92680C50EE1FC3B341F4AAF00C08EF42600C18C80E700E1FC218D00C08E",
         INIT_01 => x"54545454A6E6D0DF8E104444444462A6363439F92708C50EE1FC39F22740C50E",
         INIT_02 => x"FCBD8435FD265A20C60434B63562E762EA62A70F8462A65858585853A6E6E4E7",
         INIT_03 => x"0234A80117F12631813D273981230217F92653812A0217E2DF7F7A02171186F9",
         INIT_04 => x"E0EB02340C2904358E01170434E46AE46AE4EBE0EBE0E6103421299101172629",
         INIT_05 => x"0117E26F2402161386E2DF732C02173F86BA27FFC102355FEB2080A70527E46A",
         INIT_06 => x"2320008310062762A3E4EC0B02171286F9FCBDE4AF0130492562AC4D2930344A",
         INIT_07 => x"1780A684EB63EB62EB68011762AE750117981F03CB2F0017F3FE8E64E720C602",
         INIT_08 => x"10347120028D396532C901171486C326E4AC62AF5B0117981F53F526646A6501",
         INIT_09 => x"8D618D394AAF0229F68DF28D910017E50016F80016B301169035690017A4FE8E",
         INIT_0a => x"498D3944AF0229D58DD18D5E8D3946AF0229E08DDC8D728D3948AF0229EB8DE7",
         INIT_0b => x"8D3941A70229B18DB08D588D3942A70229BC8DBB8D6C8D3943A70229C78DC68D",
         INIT_0c => x"BF0016311FF48DB6FE8E39F726048180A651011739C4A7808A0429A68DA58D5F",
         INIT_0d => x"8DC8FE8EE12044AED78DCEFE8EB4001643A6E18DD4FE8EF42048AEEA8DC2FE8E",
         INIT_0e => x"D02042A6B38DDFFE8ED92041A6BC8DDAFE8ECF204AAEC58DBCFE8ED82046AECE",
         INIT_0f => x"B2FE8EBF8DB88DB08DA98DA18D27FF17B2FE8E900016EBFE8EC4A6AA8DE4FE8E"
      )
      port map (
         clk     => clk,
         en      => en(1),
         we      => we,
         rst     => rst,
         addr    => addr(8 downto 0),
         di      => wdata,
         do      => xdata(1)
      );

   ROM02: RAMB4_S8
      generic map (
         INIT_00 => x"3C29088D011F42290E8DCA00172D86121F4D29098DD520CE8DC78DC08D17FF17",
         INIT_01 => x"811D2530815B8D39E0AB04342829078D891F484848483229118D903561A71034",
         INIT_02 => x"3439021A39578003226681072561813937800322468112254181393080032239",
         INIT_03 => x"C602346320078B022F3981308B0F840235048D4444444402340235028D023510",
         INIT_04 => x"207F84048D0627E2DF7D00F09F6E8235F1265A518D558D2D860225E46880A608",
         INIT_05 => x"DF9FA75186EE27018584A620E08E0926018584A6E0DFBEE0DF9FA7118610343F",
         INIT_06 => x"2086008D8235018520E0B605260185E0DF9FA6E0DF9FA711860234903501A6E0",
         INIT_07 => x"84A70386E0DFBE138D903501A70235F6260885FA27028584A6E0DFBE1234498D",
         INIT_08 => x"02C6FDDFFD04E703E702A7FBDFFD0000CC30E08E39E2DFB7FF86016D84A75186",
         INIT_09 => x"20098D042420810D20608D0427FEDF7D30E08E16345986028D1B86FEDF7F01E7",
         INIT_0a => x"890027100D81382716817C0027101A815A271B81342708819635AF001784A705",
         INIT_0b => x"6D205A34275DFBDFFC8F0016792619C15CFBDFFC45260A810F270B8124270C81",
         INIT_0c => x"598114273DC1FEDFF656200000CC5820212750814CFBDFB662204A2C27FBDFB6",
         INIT_0d => x"2080FEDF7F39FDDFB70426FDDF7D39FEDF7F39FEDFB704263D81312754816E27",
         INIT_0e => x"A74C84E720C6FBDFB6168D0000CC1B20E12218C120C0FDDF7FFDDFF6ED224F81",
         INIT_0f => x"C15C4FF02650814CFBDFFC3903E702A7FBDFFDFCDFF64F39FEDF7FF726508102"
      )
      port map (
         clk     => clk,
         en      => en(2),
         we      => we,
         rst     => rst,
         addr    => addr(8 downto 0),
         di      => wdata,
         do      => xdata(2)
      );

   ROM03: RAMB4_S8
      generic map (
         INIT_00 => x"2650C15C84A702E7FBDFF72086FBDFF604E75F012519C15C04E6E78D5AEA2619",
         INIT_01 => x"FB0274FB0139FEDFF702E7FBDFF75FE4205F03E7FCDFF7082719C15CFCDFF6F4",
         INIT_02 => x"505EFA4CA5F847FDF8455CF94248FB1953FB183DFB1531FB105EFB047FFB0369",
         INIT_03 => x"94F9A7F8A7F8A7F8A7F894F992FC55D5F94488F958F1F853EDFB52A8F84DBCFA",
         INIT_04 => x"20205353455820524F4620362E312047554239305359530000000A0DFFFFFFFF",
         INIT_05 => x"43502020043D5053202004202D20043F54414857043E040000000A0D4B04202D",
         INIT_06 => x"20043D412020043D50442020043D58492020043D59492020043D53552020043D",
         INIT_07 => x"0000000000000000000004315343565A4E4948464504203A43432020043D4220",
         INIT_08 => x"300B2784AC1084AF1084EEAA558E10A0D08E84A7F086FB264A80A70F86F0FF8E",
         INIT_09 => x"2DA7D0DF8E10C0DFCE10FDFFB74444444443101F84EFD620ED26A0F08C00F089",
         INIT_0a => x"1084AF10AA558E1084EE2227A0F08C00F08930FB2A4AA66F0C862FA7F0862E6F",
         INIT_0b => x"2EA7D0DF8E10F186D520A5A70F88891F44444444101FD0DF8E1084EFE92684AC",
         INIT_0c => x"8EF32D0C814C80E7A66F0427A6E6211F4F2CE7A66F1420F92A4A0526A6E60C86",
         INIT_0d => x"9F6EC6DF9F6EC4DF9F6EC0DF9F6E62F816E2DFF753F9265A80A7A0A610C6F0FF",
         INIT_0e => x"0822CEDFBC8B300F27FFFF8CCCDFBE49584F4AAF80E64AAE431FCADF9F6EC8DF",
         INIT_0f => x"00FFB2FFC2FFBEFFBAFFB6FFC6FFB2FFC2DF9F6E42EE1F37F16E44AEC4EC1034"
      )
      port map (
         clk     => clk,
         en      => en(3),
         we      => we,
         rst     => rst,
         addr    => addr(8 downto 0),
         di      => wdata,
         do      => xdata(3)
      );

   rom_glue: process (cs, rw, addr, xdata)
   begin
      en <= (others=>'0');
      case addr(10 downto 9) is
      when "00" =>
         en(0)  <= cs;
         rdata  <= xdata(0);
      when "01" =>
         en(1)  <= cs;
         rdata  <= xdata(1);
      when "10" =>
         en(2)  <= cs;
         rdata  <= xdata(2);
      when "11" =>
         en(3)  <= cs;
         rdata  <= xdata(3);
      when others =>
         null;
      end case;
      we <= not rw;
   end process;
end architecture rtl;

