    INIT_00 => x"F9E8FAB4FBDDFB0CFABAFA15FBCEFAA5FAE9F7A5F7FEFA7BFADFF8F0F85EF17E",
    INIT_01 => x"00000200000000000000003000F3FB1F000000000003037AEA0FFDC1ED63FA61",
    INIT_02 => x"003B00003B00003B00003B00000A000000000000000003000003000000000000",
    INIT_03 => x"20375449584504020000846E0635011F45545543455845070200003B00003B00",
    INIT_04 => x"0000B16E20370227063500008310455552542D4E4F2D544958450C040000B16E",
    INIT_05 => x"4404040000B16E2037022606350000831045534C41462D4E4F2D544958450D04",
    INIT_06 => x"6E101F063410352035203653454F444F4406040000B16E10362037211F455649",
    INIT_07 => x"36EEC0BD3A4F44030400007EC03DCDD5C0BDEEC0BD52454F444F4406040000B1",
    INIT_08 => x"05040000B16E101F06341035EEC0BD4554414552434F440804BEC0B16E203520",
    INIT_09 => x"341035EEC0BD4E4F43434F4406040000B16E101F06341035EEC0BD5241564F44",
    INIT_0a => x"4F440504E4C0B16E84EC06341035EEC0BD4E4F434F440504F8C0B16E1D84E606",
    INIT_0b => x"EC06341035EEC0BD524156494F4406045DC1B16E84EC06341035EEC0BD4C4156",
    INIT_0c => x"41564F440604CEC0B16E94EC06341035EEC0BD4C4156494F4406041FC1B16E84",
    INIT_0d => x"1D5A012702845F00B0B606343F54494D45050285C0B16EE1E34958EEC0BD5352",
    INIT_0e => x"552106060000B16E063501E7FA27028484A600B08E54494D4528050486C1B16E",
    INIT_0f => x"2701845F00B0B606343F59454B04020000B16E063584A7558600B08E54524153",
    INIT_10 => x"070468C0B16E4F01E6FA2701C484E600B08E063459454B0302F2C1B16E1D5A01",
    INIT_11 => x"C4AE063424454E494C4E49070479C0B16EC4AF81ECC4AE063423454E494C4E49",
    INIT_12 => x"C4AF853080E6C4AE063424454E494C4E492F08040000B16EC4AF3A10344F80E6",
    INIT_13 => x"3500008310292846490404A1C0B16EA4AE1029284F544F47060434C2B16E0635",
    INIT_14 => x"052706350000831029284F52455A4649080476C2B16E2231B16EA4AE10052606",
    INIT_15 => x"A0E6063429432803040000B16EA1EC0634292802040000B16E2231B16EA4AE10",
    INIT_16 => x"84E3A1AE29284F542B050467C2B16E063584EDA1AE29284F540404B8C2B16E1D",
    INIT_17 => x"C2B16E063584ED0100C384EC0634A1AE292852434E4906041FC2B16E063584ED",
    INIT_18 => x"05040000B16E063510368B300636E1A30080CC011F1036A1AE29284F440404C6",
    INIT_19 => x"EC06342928504F4F4C060402C3B16EA4AE1006356232DD26E4A31029284F443F",
    INIT_1a => x"504F4F4C2B070408C2B16E063546332231B16EA4AE100635C4ED09290100C3C4",
    INIT_1b => x"33504F4F4C4E550602D6C2B16E20374433455641454C0502ACC2DE20C4E32928",
    INIT_1c => x"0493C3B16E48A346EC06344A01029BC1B16E42A3C4EC0634490102AEC1B16E46",
    INIT_1d => x"54060449C1250090C1BD47534D504F54060469C3230090C1BD434F56504F5406",
    INIT_1e => x"444C480304BEC3290090C1BD41464E504F54060408C1270090C1BD584650504F",
    INIT_1f => x"0090C1BD23534303041FC32D0090C1BD545845544E4F4307044DC22B0090C1BD",
    INIT_20 => x"04E9C2330090C1BD45444F4D0404E8C3310090C1BD322D2347534D0604DDC12F",
    INIT_21 => x"03048FC2370090C1BD53454D495423060478C3350090C1BD4E4F495443455307",
    INIT_22 => x"0090C1BD45524548540504A0C33B0090C1BD424902045AC3390090C1BD424923",
    INIT_23 => x"4D4948050636C3410090C1BD5245560306CDC33F0090C1BD524F48030633C13D",
    INIT_24 => x"C3470090C1BD3F544F44040656C4450090C1BD4B4F020604C4430090C1BD4D45",
    INIT_25 => x"BD4E493E030270C44B007BC1BD445257030420C4490090C1BD455245480402AF",
    INIT_26 => x"C453007BC1BD4554415453050230C451007BC1BD45534142040271C14F007BC1",
    INIT_27 => x"2705068AC458007BC1BD3249575327050613C455007BC1BD334957532705064B",
    INIT_28 => x"C1BD4957532704060CC55E007BC1BD515249270406E2C45B007BC1BD51524946",
    INIT_29 => x"C100C052C1BD4E494749524F06023FC464007BC1BD494D4E27040619C561007B",
    INIT_2a => x"C37F3DC1BD544E45525255430704F0C4753DC1BD4B43415453444E49460904C5",
    INIT_2b => x"0152C1BD3052020495C47E0152C1BD3053020433C5800052C1BD4249540304DC",
    INIT_2c => x"070484C5FC0252C1BD305343030486C3000252C1BD465542594C460604A2C4FE",
    INIT_2d => x"BD455552540402BBC4023DC1BD4C4C454304066EC57E3DC1BD455A4953424954",
    INIT_2e => x"4C430704F8C3203DC1BD4C4202029FC5003DC1BD45534C41460502C7C4FF3DC1",
    INIT_2f => x"0493C5B16EFE01CE522D5241454C430704AEC5B16E06357E01CE10532D524145",
    INIT_30 => x"35011F21430202DDC5B16E301F06344050520304BAC5B16E401F063440505303",
    INIT_31 => x"0635011F21320202C6C5B16E063584ED0635011F21010253C5B16E063584E706",
    INIT_32 => x"0306D4C4B16E063584ED84E30635011F212B0202FEC4B16E063584ED063581ED",
    INIT_33 => x"3584ED0100C384EC011F212B31030600C6B16E063584E784EB0635011F212B43",
    INIT_34 => x"32020279C5B16E84EC011F40010242C5B16E4F84E6011F40430202F0C5B16E06",
    INIT_35 => x"060DC6B16E10344F80E6011F544E554F43050272C6B16E103484AE81EC011F40",
    INIT_36 => x"3706343E5202027CC4B16E06350636523E0202D3C5B16E103481EC011F2B4002",
    INIT_37 => x"37063706343E52320302CEC6B16E0635063610361035523E3203029EC6B16E06",
    INIT_38 => x"C4EC103442AE06344052320302C0C6B16EC4EC063440520202E6C6B16E103410",
    INIT_39 => x"0225C7B16E4433504F52445232060608C7B16E4233504F5244520506DAC6B16E",
    INIT_3a => x"04024FC7B16E10340634E4AE505544320402F7C6B16E06356232504F52443205",
    INIT_3b => x"C7B16E66EC063466EC06345245564F3205025FC7B16E10346432103550494E32",
    INIT_3c => x"5432050264C4B16E62AF62EC1037E4ED64AF64ECE4AE06365041575332050240",
    INIT_3d => x"C088C7FBC688C7EAC6FFC0BD544F5232040232C77EC075C788C7FFC0BD4B4355",
    INIT_3e => x"C6B16E0635504F5244040293C6B16E06340227000083105055443F0402AEC67E",
    INIT_3f => x"504157530402AFC4B16E62EC06345245564F040286C6B16E0634505544030239",
