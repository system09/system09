--
-- KBUG9S

-- 4 September 2004

--

library IEEE;

  use IEEE.STD_LOGIC_1164.ALL;

  use IEEE.STD_LOGIC_ARITH.ALL;

library unisim;
	
  use unisim.vcomponents.all;



entity mon_rom is
    
  Port (

       clk   : in  std_logic;

       rst   : in  std_logic;

       cs    : in  std_logic;

       rw    : in  std_logic;

       addr  : in  std_logic_vector (10 downto 0);

       rdata : out std_logic_vector (7 downto 0);

       wdata : in  std_logic_vector (7 downto 0)

    );

end mon_rom;



architecture rtl of mon_rom is

   



signal we : std_logic;

signal dp : std_logic;



begin


  ROM : RAMB16_S9
    generic map (
 
 
    INIT_00 => x"A780A610C6C0DF8E105BFE8E6BFA6FFC73FC7FFCAEFCA0FC8BFC91FC61F814F8",
    INIT_01 => x"17431FE4A7D0866AAFDD8C30FB265AE26F0CC6F10117E0DFBF20E08EF9265AA0",
    INIT_02 => x"041783FE8EE50317F62A5A19048B0327856D0DC64FD0DF8E3704176BFE8E8604",
    INIT_03 => x"17408B981F3304175E86092C2081891FF1270D817F842704170804178AFE8E1E",
    INIT_04 => x"20E003178CFE8EF5265BFE8C02300F2780E125FE8E20C0022F60C12704172C04",
    INIT_05 => x"92FE8EF10217E90217E10217D90217D10217C1031792FE8E3B341FBC2094ADC0",
    INIT_06 => x"AD0217394AAF0229170317D70317E70217080316010317FA0217F30217AC0317",
    INIT_07 => x"17AD0317A702173946AF0229FB0217BB0317C002173948AF0229090317C90317",
    INIT_08 => x"0229E10217910317B502173943A70229EF02179F03178E02173944AF0229ED02",
    INIT_09 => x"C4A7808A0429C50217750317A302173941A70229D302178303179D02173942A7",
    INIT_0a => x"02174E0317E50217A4A6560317E50217211F21031792FE8E121F2D29AB021739",
    INIT_0b => x"173F862F03170827A4A1A4A7390F260D8117275E81DD271881E127088111289E",
    INIT_0c => x"24E1AC203406294B021705201F30C0DF8E321FF50117BE203F31C22021312C03",
    INIT_0d => x"8E10343962320327E802170527E4AC011FF0C4201F0634F0C41000C3101F3901",
    INIT_0e => x"80A610C6E1AED00217F5265AD802176F021780A610C66E0217E4AEAA021792FE",
    INIT_0f => x"FF8E10341A24C0DF8C1E29FA0117BF20EE265AC102172E8602237E8104252081",
    INIT_10 => x"8E109002163F869302173984A73F86A4AFA0A709273F8184A60F271035558DFF",
    INIT_11 => x"21AE23FE166DFE17068D4AAF0427268D1F304AAE431F39FB265A188D08C6E3DF",
    INIT_12 => x"A0A608C6E3DF8E1039A0A7A0A7A0A7FF8684A7A4A604263F8184A60A24C0DF8C",
    INIT_13 => x"E6E4E754545454A6E6D0DF8E104444444462A63634393D3139F7265A0427A1AC",
    INIT_14 => x"DFBF00E08E8435FD265A20C60434B63562E762EA62A70F8462A65858585853A6",
    INIT_15 => x"0117F126318149273981D00117F9265381D70117E2DF7F0502171186C8FCBDE0",
    INIT_16 => x"340C2904352401170434E46AE46AE4EBE0EBE0E610342129270117262902343E",
    INIT_17 => x"00E08EB101173F86E0DFBF20E08EBA27FFC102355FEB2080A70527E46AE0EB02",
    INIT_18 => x"304F2562AC53293034CD0017E26F39E0DFBF20E08EA301171386E2DF73E0DFBF",
    INIT_19 => x"E720C6022320008310062762A3E4EC7D01171286C8FCBDE0DFBF00E08EE4AF01",
    INIT_1a => x"646AE2001780A684EB63EB62EBE5001762AEF20017981F03CB280117FAFE8E64",
    INIT_1b => x"DFBF20E08E65323501171486E0DFBF00E08EC326E4AC62AFD80017981F53F526",
    INIT_1c => x"43A6E10017DBFE8EA0001648AEEC0017C9FE8EAB0016311FF70017BDFE8E39E0",
    INIT_1d => x"AEC00017C3FE8E7F001646AECB0017CFFE8E8A001644AED60017D5FE8E9D0016",
    INIT_1e => x"8EC4A6A20017EBFE8E692042A6AC0017E6FE8E732041A6B60017E1FE8E75204A",
    INIT_1f => x"8D903561A710343C29088D011F42290E8DBF00172D86121F4D29098D7220F2FE",
    INIT_20 => x"81393080032239811D253081728D39E0AB04342829078D891F48484848322911",
    INIT_21 => x"0235028D0235103439021A395780032266810725618139378003224681122541",
    INIT_22 => x"0225E46880A608C602345820078B022F3981308B0F840235048D444444440234",
    INIT_23 => x"A62F8D391035058D84FE8E10340C20028D00F09F6E8235F1265A468D4A8D2D86",
    INIT_24 => x"903501A6FA27018584A6E0DFBE10341D207F84048D0627E2DF7D39F826048180",
    INIT_25 => x"028584A69235458D042620E08CE0DFBE12342086008D82350185E0DF9FA60234",
    INIT_26 => x"39012720E08CE2DFB7FF86016D84A7118684A70386E0DFBE903501A70235FA27",
    INIT_27 => x"345986028D1B86FEDF7F01E702C6FDDFFD04E703E702A7FBDFFD0000CC30E08E",
    INIT_28 => x"271008819635C5001784A70520098D042420810D20748D0427FEDF7D30E08E16",
    INIT_29 => x"2C0027100C81990027100D814500271016818E0027101A816C0027101B814100",
    INIT_2a => x"5A3C0027105DFBDFFC9900168300261019C15CFBDFFC51260A81110027100B81",
    INIT_2b => x"F65800160000CC5B00162500271050814CFBDFB66800164A3327FBDFB6740016",
    INIT_2c => x"26FDDF7D39FEDF7F39FEDFB704263D81312754816E002710598116273DC1FEDF",
    INIT_2d => x"8D0000CC1B20E12218C120C0FDDF7FFDDFF6ED224F812080FEDF7F39FDDFB704",
    INIT_2e => x"FC3903E702A7FBDFFDFCDFF64F39FEDF7FF726508102A74C84E720C6FBDFB616",
    INIT_2f => x"F72086FBDFF604E75F012519C15C04E6E78D5AEA2619C15C4FF02650814CFBDF",
    INIT_30 => x"E7FBDFF75FE4205F03E7FCDFF7082719C15CFCDFF6F42650C15C84A702E7FBDF",
    INIT_31 => x"F2F942EBF819F9F818DDF815CFF81007F90431F90315F90223F90139FEDFF702",
    INIT_32 => x"F8A7F82AFA6BFC551EFA588AF953A8F85241F94D12FB509BFA4CA5F84796F945",
    INIT_33 => x"20312E312047554239305359530000000A0D000000FFFFFFFF2AFAA7F8A7F8A7",
    INIT_34 => x"202C042053534150202C04202D20043F54414857043E040000000A0D4B04202D",
    INIT_35 => x"532020303132333435363704203E3D2004203A524F525245204E492053544942",
    INIT_36 => x"3D50442020043D58492020043D59492020043D53552020043D43502020043D50",
    INIT_37 => x"00000004315343565A4E4948464504203A43432020043D422020043D41202004",
    INIT_38 => x"300B2784AC1084AF1084EEAA558E10A0D08E84A7F086FB264A80A70F86F0FF8E",
    INIT_39 => x"2DA7D0DF8E10C0DFCE10FDFFB74444444443101F84EFD620ED26A0F08C00F089",
    INIT_3a => x"1084AF10AA558E1084EE2227A0F08C00F08930FB2A4AA66F0C862FA7F0862E6F",
    INIT_3b => x"2EA7D0DF8E10F186D520A5A70F88891F44444444101FD0DF8E1084EFE92684AC",
    INIT_3c => x"8EF32D0C814C80E7A66F0427A6E6211F4F2CE7A66F1420F92A4A0526A6E60C86",
    INIT_3d => x"9F6EC6DF9F6EC4DF9F6EC0DF9F6E62F816E2DFF753F9265A80A7A0A610C6F0FF",
    INIT_3e => x"0822CEDFBC8B300F27FFFF8CCCDFBE49584F4AAF80E64AAE431FCADF9F6EC8DF",
    INIT_3f => x"00FFB2FFC2FFBEFFBAFFB6FFC6FFB2FFC2DF9F6E42EE1F37F16E44AEC4EC1034"
   )


    port map (

	  do     => rdata,

	  dop(0) => dp,

	  addr   => addr,

	  clk    => clk,

	  di     => wdata,

	  dip(0) => dp,

	  en     => cs,

	  ssr    => rst,

	  we     => we

	);



my_mon : process ( rw )

begin

	 we    <= not rw;

end process;



end architecture rtl;

