    INIT_00 => x"ACFC8E1001E07D00E0B7118600E0B70386FA2612121F3000008E20F6CE10321A",
    INIT_01 => x"2AF6B72BF6B72EF6FD0000CC22F6F723F6B710F6CCFA265A81AF1008C600F08E",
    INIT_02 => x"34D1FD7E30F6B7FA862DF6B7828621F6B720F6B724F6FD26F6FD28F6FD2CF6B7",
    INIT_03 => x"FCBD02349035011A903501E0B64FF227018400E0B60D271F308EFCBD00008E10",
    INIT_04 => x"6D20393038363F0100000000008005394C4F3901E0B70235F627028400E0B68E",
    INIT_05 => x"02352AF6B702352BF6B702352DF6B7023520F6B700302E315620726F74696E6F",
    INIT_06 => x"20F6B6103524F6F725F6B7063526F6F727F6B7063528F6F729F6B706352CF6B7",
    INIT_07 => x"25F781F4255FFCBD30F68E20F6CE1037FE7E2EF6F72FF6B7101F1F3002260181",
    INIT_08 => x"FCBDF6265A80A7D8255FFCBD891F0C27008180A7E5228081E9255FFCBD80A7F0",
    INIT_09 => x"812527FD812627FE814227FF8180E680A630F68EC526E0ABB4FEBD0234CE255F",
    INIT_0a => x"FE7E018630F6B7F0861F27F7812027F8812127F9812227FA812327FB812427FC",
    INIT_0b => x"31F68E1091FC8E84FE7E79FE7E4BFE7EF8FD7EE6FD7ED1FD7EA5FD7E8EFD7E92",
    INIT_0c => x"5A80A7A0A6072731F6F703E6021F01E602A69CFE7EF9265AA0A780A6A0E71BC6",
    INIT_0d => x"A63435F9265AA0A780A63434142703C031F6F6021F80A680E680A69CFE7EF926",
    INIT_0e => x"80A7A0A680E731F68E10C620F68E1092FE7E018602200086F7265A0726A0A180",
    INIT_0f => x"041F22F6F623F6B692FE7E4FF9265AA0A780A620F68E100B275D9CFE7EF9265A",
