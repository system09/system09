--===========================================================================--
--                                                                           --
--    Synthesizable Character Generator using Xilinx RAMB16_S9 Block RAM     --
--                                                                           --
--===========================================================================--
--
--  File name      : char_rom2k_b16.vhd
--
--  Entity name    : char_rom
--
--  Purpose        : Implements a character generator ROM
--                   using one Xilinx RAMB16_S9 Block RAM
--                   Used by vdu8.vhd in the System09 SoC
--
--  Dependencies   : ieee.std_logic_1164
--                   ieee.std_logic_arith
--
--  Uses           : RAMB16_S9 (Xilinx 16KBit Block RAM)
--
--  Author         : John E. Kent
--
--  Email          : dilbert57@opencores.org      
--
--  Web            : http://opencores.org/project,system09
--
--  Description    : Characters are 7 pixels x 11 rows x 128 characters
--                   Stored as 8 bits x 16 locations x 128 characters
--
--  Copyright (C) 2003 - 2010 John Kent
--
--  This program is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
--===========================================================================--
--                                                                           --
--                              Revision  History                            --
--                                                                           --
--===========================================================================--
--
-- Version Date        Author     Changes
--
-- 0.1     2004-10-18  John Kent  Initial relaease
--
-- 0.2     2010-06-17  John Kent  Updated header and description and added GPL
--     

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
library unisim;
	use unisim.vcomponents.all;

entity char_rom is
    Port (
       clk      : in  std_logic;
       rst      : in  std_logic;
       cs       : in  std_logic;
       addr     : in  std_logic_vector (10 downto 0);
       rw       : in  std_logic;
       data_in  : in  std_logic_vector (7 downto 0);
       data_out : out std_logic_vector (7 downto 0)
    );
end char_rom;

architecture rtl of char_rom is


signal we : std_logic;
signal dp : std_logic;

begin

  ROM : RAMB16_S9
    generic map (
    INIT_00 => x"000000000009090F09090038043840380000000000070404040400444C546444",
    INIT_01 => x"0000000000110A040A110078407040780000000000110A040A11003804384038",
    INIT_02 => x"00000000000D1215110E0078407040780000000000040404041F007840704078",
    INIT_03 => x"00000000000F080808080070487048700000000000090A0C0A09004878484830",
    INIT_04 => x"0000000000040404041F0044447C444400000000000E010E100E007048704870",
    INIT_05 => x"0000000000040404041F001028444444000000000010101E101F007C40404040",
    INIT_06 => x"000000000011111E111E003C4040403C000000000008080E080F004040704078",
    INIT_07 => x"0000000000070202020700380438403800000000000E1111110E003804384038",
    INIT_08 => x"0000000000070202060200704848487000000000000F080E080F007048484870",
    INIT_09 => x"00000000000E0107020F00704848487000000000000F08060907007048484870",
    INIT_0a => x"0000000000090A0C0A0900444C546444000000000001010F0909007048484870",
    INIT_0b => x"00000000000E090E090E00784070407800000000001113151911003804384038",
    INIT_0c => x"00000000001111151B1100784070407800000000001113151911003840404038",
    INIT_0d => x"00000000000E1010100E00784070407800000000000E090E090E003804384038",
    INIT_0e => x"00000000000E010E100E00384858403800000000000E010E100E004040704078",
    INIT_0f => x"00000000000E010E100E00304848484800000000000E010E100E004850704870",
    INIT_10 => x"0000000000080800000808080808080800000000000000000000000000000000",
    INIT_11 => x"00000000002424247E2424247E24242400000000000000000000000012121212",
    INIT_12 => x"000000000043434020100804020161610000000000083E4909093E4848493E08",
    INIT_13 => x"0000000000000000000000002010080C00000000003D42444444384444444438",
    INIT_14 => x"0000000000201008040404040408102000000000000204081010101010080402",
    INIT_15 => x"000000000000000808087F0808080000000000000000004122147F1422410000",
    INIT_16 => x"000000000000000000007F000000000000004020101818000000000000000000",
    INIT_17 => x"0000000000404040201008040201010100000000001818000000000000000000",
    INIT_18 => x"00000000003E0808080808080828180800000000000814224141414141221408",
    INIT_19 => x"00000000003E410101010E010101413E00000000007F4020100804020141423C",
    INIT_1a => x"00000000003E410101615E404040407F000000000002020202027F22120A0602",
    INIT_1b => x"0000000000404020100804020101017F00000000001E214141615E404040211E",
    INIT_1c => x"00000000003C420101013D434141423C00000000003E414141413E414141413E",
    INIT_1d => x"0000004020101818180000001818180000000000000018181800000018181800",
    INIT_1e => x"0000000000000000007F00007F00000000000000000102040810201008040201",
    INIT_1f => x"0000000000080800080808060101413E00000000004020100804020408102040",
    INIT_20 => x"000000000041414141417F414122140800000000001C224140404E494541221C",
    INIT_21 => x"00000000001E2141404040404041211E00000000007E212121213E212121217E",
    INIT_22 => x"00000000007F404040407C404040407F00000000007C2221212121212121227C",
    INIT_23 => x"00000000001E2141414147404040211E000000000040404040407C404040407F",
    INIT_24 => x"00000000003E0808080808080808083E000000000041414141417F4141414141",
    INIT_25 => x"0000000000414244485060504844424100000000003C42020202020202020207",
    INIT_26 => x"0000000000414141414141494955634100000000007F40404040404040404040",
    INIT_27 => x"00000000003E4141414141414141413E00000000004141414345494951614141", -- 
    INIT_28 => x"00000000003D4245494141414141413E000000000040404040407E414141417E", -- P Q
    INIT_29 => x"00000000003E410101013E404040413E000000000041424448507E414141417E", -- R S
    INIT_2a => x"00000000003E414141414141414141410000000000080808080808080808087F", -- T U
    INIT_2b => x"0000000000222255554949414141414100000000000808141414222222414141", -- V W
    INIT_2c => x"0000000000080808080808142241414100000000004141412214081422414141", -- X Y
    INIT_2d => x"00000000001E1010101010101010101E00000000007F4040201008040201017F", -- Z [
    INIT_2e => x"00000000003C0404040404040404043C00000000000101010204081020404040", -- \ ]
    INIT_2f => x"00000000007F0000000000000000000000000000000000000000000041221408", -- _ ^
    INIT_30 => x"00000000003F41413F01013E0000000000000000000000000000000002040818", -- ` a
    INIT_31 => x"00000000001E21404040211E0000000000000000005E61616141615E40404040", -- b c
    INIT_32 => x"00000000003E40407F41413E0000000000000000003D43414141433D01010101", -- d e
    INIT_33 => x"00003C4202023E424242423D0100000000000000001010101010107C1010110E", -- f g
    INIT_34 => x"00000000003E0808080808180000080800000000004141414141615E40404040", -- h i
    INIT_35 => x"0000000000414448704844414040404000003C42020202020202020200000202", -- j k
    INIT_36 => x"0000000000414141494955220000000000000000001C08080808080808080818", -- l m
    INIT_37 => x"00000000003E41414141413E0000000000000000004141414141615E00000000", -- n o
    INIT_38 => x"0000010101013D434343433D000000000000404040405E616161615E00000000", -- p q
    INIT_39 => x"00000000003E01013E40403E0000000000000000002020202020314E00000000", -- r s
    INIT_3a => x"00000000003D4242424242420000000000000000000C12101010107C10101010", -- t u
    INIT_3b => x"0000000000225549494141410000000000000000000814142222414100000000", -- v w
    INIT_3c => x"00003C4202023A46424242420000000000000000004122140814224100000000", -- x y
    INIT_3d => x"0000000000070808081020100808080700000000007F20100804027F00000000", -- z {
    INIT_3e => x"0000000000700808080402040808087000000000000808080808000808080808", -- | }
    INIT_3f => x"0000000000492249224922492249224900000000000000000000000000464931"  -- ~ del
    )

    port map (
	  do    => data_out,
	  dop(0)=> dp,
	  addr  => addr,
	  clk   => clk,
     di    => data_in,
	  dip(0)=> dp,
	  en    => cs,
	  ssr   => rst,
	  we    => we
	);

my_char_rom : process ( rw )
begin
	 we    <= not rw;
end process;

end architecture rtl;

