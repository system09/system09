    INIT_00 => x"C725D87BC2D4C88900AFC2E6C737C98F00AFC2E6C7FFC0BD44455845444E4907",
    INIT_01 => x"C2D4C88F00AFC2E6C77EC066D7DBC737D87BC2D4C88D00AFC2E6C77EC09ED7DB",
    INIT_02 => x"C989C6FFC0BD44454D4D4905043AD77EC0FDCCDBC77EC0E8CCFDCCDBC74BD87B",
    INIT_03 => x"D5C0BDEEC0BD5845534F44050468D67EC0FDCC7EC0E8CC6DD87BC2B8D646CEB9",
    INIT_04 => x"7EC0A0D6E8CC95C6D5C0BDEEC0BD324957534F44060487D57EC0A0D6FDCC89C6",
    INIT_05 => x"ABD57EC0A0D6FDCCFDCC89C6B8D618C4D5C0BDEEC0BD494157434F44060419D4",
    INIT_06 => x"7EC05AD8DBC7E0D87BC2D4C800BCC2E6C7A0D618C4FFC0BD5244414E45470604",
    INIT_07 => x"DBC706D97BC2D4C820BCC2E6C77EC0FDCCDBC7DBC7F3D87BC2D4C810BCC2E6C7",
    INIT_08 => x"04A3D87EC0B8D67EC0E8CCDBC7DBC719D97BC2D4C830BCC2E6C77EC008D8DBC7",
    INIT_09 => x"BD59444C4F44050480D67EC0C8D8FDCC40D7B4C6D5C0BDEEC0BD47454E4F4405",
    INIT_0a => x"89C6D5C0BDEEC0BD4758454F44050420D97EC0C8D8E8CC40D7C3C6D5C0BDEEC0",
    INIT_0b => x"D5C0BDEEC0BD41454C4F44050439D97EC0A0D6FDCCD7C96EC904BCC200C8FDCC",
    INIT_0c => x"BDEEC0BD5145424F44050474D97EC0A0D608D8FDCC89C6B8D6E0C920BCC218C4",
    INIT_0d => x"C0FDCCFDCC00C8C1D97BC286D6E6C7A0D6E0C9D7C902BCC2A7C400C889C6D5C0",
    INIT_0e => x"BDEEC0BD4152424F44050496D97EC0E8CCE0C902BCC2FDCC00C8FDCC10BCC27E",
    INIT_0f => x"CCFDCCA4C900C803DA7BC286D6E6C7A0D6E0C9D7C902BCC2A7C400C895C6D5C0",
    INIT_10 => x"C0D0D689C6D5C0BDEEC0BD292D4F44040499D57EC0E8CCB9C9FDCC00C87EC0FD",
    INIT_11 => x"52534C0308F3D6004329D9BD4D4F43030854D8004029D9BD47454E030860D77E",
    INIT_12 => x"0830DA004729D9BD52534103084BD6004629D9BD524F52030881D1004429D9BD",
    INIT_13 => x"4929D9BD4C4F52030810DA004829D9BD4C534C03088BD8004829D9BD4C534103",
    INIT_14 => x"545354030874D8004C29D9BD434E49030897D7004A29D9BD434544030852D900",
    INIT_15 => x"0812D5004F29D9BD524C430308C1D8004E29D9BD504D4A030878DA004D29D9BD",
    INIT_16 => x"BD414342530408CDDA018129D9BD41504D430408C0DA018029D9BD4142555304",
    INIT_17 => x"9CDA018429D9BD41444E41040890DA028329D9BD444255530408B4DA018229D9",
    INIT_18 => x"D9BD415453030800D8018629D9BD41444C0308D6D9018529D9BD415449420408",
    INIT_19 => x"08DADA018929D9BD414344410408F4DA018829D9BD41524F450408C7D6008729",
    INIT_1a => x"D9BD58504D4304084CDB018B29D9BD41444441040833DB018A29D9BD41524F03",
    INIT_1b => x"5303082BD6028E29D9BD58444C030801DB008D29D9BD52534A03080EDB028C29",
    INIT_1c => x"C129D9BD42504D4304088ADB01C029D9BD42425553040826DB008F29D9BD5854",
    INIT_1d => x"41040860DA02C329D9BD44444441040854DA01C229D9BD42434253040897DB01",
    INIT_1e => x"C629D9BD42444C03083CDA01C529D9BD425449420408A8DA01C429D9BD42444E",
    INIT_1f => x"44410408BEDB01C829D9BD42524F45040840DB00C729D9BD4254530308E7DA01",
    INIT_20 => x"01CB29D9BD424444410408FDDB01CA29D9BD42524F0308A4DB01C929D9BD4243",
    INIT_21 => x"BD55444C030848DA00CD29D9BD44545303080ADC02CC29D9BD44444C03086CDA",
    INIT_22 => x"F0DB02831042D9BD44504D430408E4DB00CF29D9BD555453030816DC02CE29D9",
    INIT_23 => x"59545303081ADB028E1042D9BD59444C030866DB028C1042D9BD59504D430408",
    INIT_24 => x"00CF1042D9BD5354530308B1DB02CE1042D9BD53444C0308CBDB008F1042D9BD",
    INIT_25 => x"040824DA028C1142D9BD53504D43040847DC02831142D9BD55504D43040896DC",
    INIT_26 => x"327DD9BD5341454C04083BDC317DD9BD5941454C040884DA307DD9BD5841454C",
    INIT_27 => x"D9BD5246540308BFDC1E5BD9BD47584503082FDC337DD9BD5541454C040889DC",
    INIT_28 => x"4141440308D7DC137DD8BD434E59530408B1DC127DD8BD504F4E03086FDC1F5B",
    INIT_29 => x"424103087CDC397DD8BD535452030823DC1D7DD8BD58455303087EDB197DD8BD",
    INIT_2a => x"5303083DDD3D7DD8BD4C554D0308A3DC3B7DD8BD4954520308FADC3A7DD8BD58",
    INIT_2b => x"CBDC437DD8BD414D4F43040861DC407DD8BD4147454E040848DD3F7DD8BD4957",
    INIT_2c => x"D8BD41525341040859DB467DD8BD41524F52040872DB447DD8BD4152534C0408",
    INIT_2d => x"4F5204088DDD487DD8BD414C534C040881DD487DD8BD414C5341040899DD477D",
    INIT_2e => x"C9DD4C7DD8BD41434E49040853DC4A7DD8BD414345440408E3DC497DD8BD414C",
    INIT_2f => x"D8BD4247454E04081CDD4F7DD8BD41524C43040875DD4D7DD8BD415453540408",
    INIT_30 => x"4F520408E1DD547DD8BD4252534C040832DD537DD8BD424D4F430408EFDC507D",
    INIT_31 => x"11DE587DD8BD424C5341040829DE577DD8BD42525341040810DD567DD8BD4252",
    INIT_32 => x"D8BD424345440408BDDD597DD8BD424C4F5204081DDE587DD8BD424C534C0408",
    INIT_33 => x"4C43040805DE5D7DD8BD42545354040859DE5C7DD8BD42434E4904085EDD5A7D",
    INIT_34 => x"3F1195D8BD33495753040835DE3F1095D8BD3249575304087DDE5F7DD8BD4252",
    INIT_35 => x"48535004084DDE1CADD8BD4343444E410508A5DD1AADD8BD4343524F040853DD",
    INIT_36 => x"08D4DE36ADD8BD554853500408F9DD35ADD8BD534C55500408BCDE34ADD8BD53",
    INIT_37 => x"20DFD9BD415242030869DD3CADD8BD494157430408EDDD37ADD8BD554C555004",
    INIT_38 => x"BD4948420308F8DE219FD9BD4E5242030805DD178DDFD9BD5253420308E0DE16",
    INIT_39 => x"4F4C42030871DE249FD9BD534842030826DF239FD9BD534C42030841DE229FD9",
    INIT_3a => x"4E420308D8DB259FD9BD534342030847DF249FD9BD434342030831DF259FD9BD",
    INIT_3b => x"42030873DF289FD9BD435642030852DF279FD9BD51454203081BDF269FD9BD45",
    INIT_3c => x"03085DDF2B9FD9BD494D42030868DF2A9FD9BD4C50420308C8DE299FD9BD5356",
    INIT_3d => x"089FDF2E9FD9BD5447420308AADF2D9FD9BD544C42030889DF2C9FD9BD454742",
    INIT_3e => x"ECDE243DC1BD3F3C550308CBDF233DC1BD3F3E55030889DE2F9FD9BD454C4203",
    INIT_3f => x"10DF283DC1BD3F53560308C0DF263DC1BD3F3D0208D5DD243DC1BD3F53430308",
